magic
tech sky130A
magscale 1 2
timestamp 1766711446
<< obsli1 >>
rect 1104 2159 134596 135473
<< obsm1 >>
rect 14 1912 134766 135504
<< metal2 >>
rect 18 137058 74 137858
rect 3238 137058 3294 137858
rect 6458 137058 6514 137858
rect 9678 137058 9734 137858
rect 12898 137058 12954 137858
rect 16118 137058 16174 137858
rect 19338 137058 19394 137858
rect 21914 137058 21970 137858
rect 25134 137058 25190 137858
rect 28354 137058 28410 137858
rect 31574 137058 31630 137858
rect 34794 137058 34850 137858
rect 38014 137058 38070 137858
rect 41234 137058 41290 137858
rect 44454 137058 44510 137858
rect 47674 137058 47730 137858
rect 50894 137058 50950 137858
rect 54114 137058 54170 137858
rect 57334 137058 57390 137858
rect 60554 137058 60610 137858
rect 63774 137058 63830 137858
rect 66994 137058 67050 137858
rect 70214 137058 70270 137858
rect 73434 137058 73490 137858
rect 76654 137058 76710 137858
rect 79874 137058 79930 137858
rect 83094 137058 83150 137858
rect 86314 137058 86370 137858
rect 89534 137058 89590 137858
rect 92754 137058 92810 137858
rect 95974 137058 96030 137858
rect 98550 137058 98606 137858
rect 101770 137058 101826 137858
rect 104990 137058 105046 137858
rect 108210 137058 108266 137858
rect 111430 137058 111486 137858
rect 114650 137058 114706 137858
rect 117870 137058 117926 137858
rect 121090 137058 121146 137858
rect 124310 137058 124366 137858
rect 127530 137058 127586 137858
rect 130750 137058 130806 137858
rect 133970 137058 134026 137858
rect 18 0 74 800
rect 2594 0 2650 800
rect 5814 0 5870 800
rect 9034 0 9090 800
rect 12254 0 12310 800
rect 15474 0 15530 800
rect 18694 0 18750 800
rect 21914 0 21970 800
rect 25134 0 25190 800
rect 28354 0 28410 800
rect 31574 0 31630 800
rect 34794 0 34850 800
rect 38014 0 38070 800
rect 41234 0 41290 800
rect 44454 0 44510 800
rect 47674 0 47730 800
rect 50894 0 50950 800
rect 54114 0 54170 800
rect 57334 0 57390 800
rect 60554 0 60610 800
rect 63774 0 63830 800
rect 66994 0 67050 800
rect 70214 0 70270 800
rect 73434 0 73490 800
rect 76010 0 76066 800
rect 79230 0 79286 800
rect 82450 0 82506 800
rect 85670 0 85726 800
rect 88890 0 88946 800
rect 92110 0 92166 800
rect 95330 0 95386 800
rect 98550 0 98606 800
rect 101770 0 101826 800
rect 104990 0 105046 800
rect 108210 0 108266 800
rect 111430 0 111486 800
rect 114650 0 114706 800
rect 117870 0 117926 800
rect 121090 0 121146 800
rect 124310 0 124366 800
rect 127530 0 127586 800
rect 130750 0 130806 800
rect 133970 0 134026 800
<< obsm2 >>
rect 130 137002 3182 137170
rect 3350 137002 6402 137170
rect 6570 137002 9622 137170
rect 9790 137002 12842 137170
rect 13010 137002 16062 137170
rect 16230 137002 19282 137170
rect 19450 137002 21858 137170
rect 22026 137002 25078 137170
rect 25246 137002 28298 137170
rect 28466 137002 31518 137170
rect 31686 137002 34738 137170
rect 34906 137002 37958 137170
rect 38126 137002 41178 137170
rect 41346 137002 44398 137170
rect 44566 137002 47618 137170
rect 47786 137002 50838 137170
rect 51006 137002 54058 137170
rect 54226 137002 57278 137170
rect 57446 137002 60498 137170
rect 60666 137002 63718 137170
rect 63886 137002 66938 137170
rect 67106 137002 70158 137170
rect 70326 137002 73378 137170
rect 73546 137002 76598 137170
rect 76766 137002 79818 137170
rect 79986 137002 83038 137170
rect 83206 137002 86258 137170
rect 86426 137002 89478 137170
rect 89646 137002 92698 137170
rect 92866 137002 95918 137170
rect 96086 137002 98494 137170
rect 98662 137002 101714 137170
rect 101882 137002 104934 137170
rect 105102 137002 108154 137170
rect 108322 137002 111374 137170
rect 111542 137002 114594 137170
rect 114762 137002 117814 137170
rect 117982 137002 121034 137170
rect 121202 137002 124254 137170
rect 124422 137002 127474 137170
rect 127642 137002 130694 137170
rect 130862 137002 133914 137170
rect 134082 137002 134762 137170
rect 20 856 134762 137002
rect 130 734 2538 856
rect 2706 734 5758 856
rect 5926 734 8978 856
rect 9146 734 12198 856
rect 12366 734 15418 856
rect 15586 734 18638 856
rect 18806 734 21858 856
rect 22026 734 25078 856
rect 25246 734 28298 856
rect 28466 734 31518 856
rect 31686 734 34738 856
rect 34906 734 37958 856
rect 38126 734 41178 856
rect 41346 734 44398 856
rect 44566 734 47618 856
rect 47786 734 50838 856
rect 51006 734 54058 856
rect 54226 734 57278 856
rect 57446 734 60498 856
rect 60666 734 63718 856
rect 63886 734 66938 856
rect 67106 734 70158 856
rect 70326 734 73378 856
rect 73546 734 75954 856
rect 76122 734 79174 856
rect 79342 734 82394 856
rect 82562 734 85614 856
rect 85782 734 88834 856
rect 89002 734 92054 856
rect 92222 734 95274 856
rect 95442 734 98494 856
rect 98662 734 101714 856
rect 101882 734 104934 856
rect 105102 734 108154 856
rect 108322 734 111374 856
rect 111542 734 114594 856
rect 114762 734 117814 856
rect 117982 734 121034 856
rect 121202 734 124254 856
rect 124422 734 127474 856
rect 127642 734 130694 856
rect 130862 734 133914 856
rect 134082 734 134762 856
<< metal3 >>
rect 134914 136008 135714 136128
rect 0 134648 800 134768
rect 134914 132608 135714 132728
rect 0 131248 800 131368
rect 134914 129208 135714 129328
rect 0 127848 800 127968
rect 134914 125808 135714 125928
rect 0 124448 800 124568
rect 134914 122408 135714 122528
rect 0 121048 800 121168
rect 134914 119008 135714 119128
rect 0 117648 800 117768
rect 134914 115608 135714 115728
rect 0 114248 800 114368
rect 134914 112208 135714 112328
rect 0 110848 800 110968
rect 134914 108808 135714 108928
rect 0 107448 800 107568
rect 134914 105408 135714 105528
rect 0 104048 800 104168
rect 134914 102008 135714 102128
rect 0 100648 800 100768
rect 134914 98608 135714 98728
rect 0 97248 800 97368
rect 134914 95888 135714 96008
rect 0 93848 800 93968
rect 134914 92488 135714 92608
rect 0 90448 800 90568
rect 134914 89088 135714 89208
rect 0 87048 800 87168
rect 134914 85688 135714 85808
rect 0 83648 800 83768
rect 134914 82288 135714 82408
rect 0 80248 800 80368
rect 134914 78888 135714 79008
rect 0 77528 800 77648
rect 134914 75488 135714 75608
rect 0 74128 800 74248
rect 134914 72088 135714 72208
rect 0 70728 800 70848
rect 134914 68688 135714 68808
rect 0 67328 800 67448
rect 134914 65288 135714 65408
rect 0 63928 800 64048
rect 134914 61888 135714 62008
rect 0 60528 800 60648
rect 134914 58488 135714 58608
rect 0 57128 800 57248
rect 134914 55088 135714 55208
rect 0 53728 800 53848
rect 134914 51688 135714 51808
rect 0 50328 800 50448
rect 134914 48288 135714 48408
rect 0 46928 800 47048
rect 134914 44888 135714 45008
rect 0 43528 800 43648
rect 134914 41488 135714 41608
rect 0 40128 800 40248
rect 134914 38088 135714 38208
rect 0 36728 800 36848
rect 134914 34688 135714 34808
rect 0 33328 800 33448
rect 134914 31288 135714 31408
rect 0 29928 800 30048
rect 134914 27888 135714 28008
rect 0 26528 800 26648
rect 134914 24488 135714 24608
rect 0 23128 800 23248
rect 134914 21088 135714 21208
rect 0 19728 800 19848
rect 134914 17688 135714 17808
rect 0 16328 800 16448
rect 134914 14968 135714 15088
rect 0 12928 800 13048
rect 134914 11568 135714 11688
rect 0 9528 800 9648
rect 134914 8168 135714 8288
rect 0 6128 800 6248
rect 134914 4768 135714 4888
rect 0 2728 800 2848
rect 134914 1368 135714 1488
<< obsm3 >>
rect 798 135928 134834 136101
rect 798 134848 134914 135928
rect 880 134568 134914 134848
rect 798 132808 134914 134568
rect 798 132528 134834 132808
rect 798 131448 134914 132528
rect 880 131168 134914 131448
rect 798 129408 134914 131168
rect 798 129128 134834 129408
rect 798 128048 134914 129128
rect 880 127768 134914 128048
rect 798 126008 134914 127768
rect 798 125728 134834 126008
rect 798 124648 134914 125728
rect 880 124368 134914 124648
rect 798 122608 134914 124368
rect 798 122328 134834 122608
rect 798 121248 134914 122328
rect 880 120968 134914 121248
rect 798 119208 134914 120968
rect 798 118928 134834 119208
rect 798 117848 134914 118928
rect 880 117568 134914 117848
rect 798 115808 134914 117568
rect 798 115528 134834 115808
rect 798 114448 134914 115528
rect 880 114168 134914 114448
rect 798 112408 134914 114168
rect 798 112128 134834 112408
rect 798 111048 134914 112128
rect 880 110768 134914 111048
rect 798 109008 134914 110768
rect 798 108728 134834 109008
rect 798 107648 134914 108728
rect 880 107368 134914 107648
rect 798 105608 134914 107368
rect 798 105328 134834 105608
rect 798 104248 134914 105328
rect 880 103968 134914 104248
rect 798 102208 134914 103968
rect 798 101928 134834 102208
rect 798 100848 134914 101928
rect 880 100568 134914 100848
rect 798 98808 134914 100568
rect 798 98528 134834 98808
rect 798 97448 134914 98528
rect 880 97168 134914 97448
rect 798 96088 134914 97168
rect 798 95808 134834 96088
rect 798 94048 134914 95808
rect 880 93768 134914 94048
rect 798 92688 134914 93768
rect 798 92408 134834 92688
rect 798 90648 134914 92408
rect 880 90368 134914 90648
rect 798 89288 134914 90368
rect 798 89008 134834 89288
rect 798 87248 134914 89008
rect 880 86968 134914 87248
rect 798 85888 134914 86968
rect 798 85608 134834 85888
rect 798 83848 134914 85608
rect 880 83568 134914 83848
rect 798 82488 134914 83568
rect 798 82208 134834 82488
rect 798 80448 134914 82208
rect 880 80168 134914 80448
rect 798 79088 134914 80168
rect 798 78808 134834 79088
rect 798 77728 134914 78808
rect 880 77448 134914 77728
rect 798 75688 134914 77448
rect 798 75408 134834 75688
rect 798 74328 134914 75408
rect 880 74048 134914 74328
rect 798 72288 134914 74048
rect 798 72008 134834 72288
rect 798 70928 134914 72008
rect 880 70648 134914 70928
rect 798 68888 134914 70648
rect 798 68608 134834 68888
rect 798 67528 134914 68608
rect 880 67248 134914 67528
rect 798 65488 134914 67248
rect 798 65208 134834 65488
rect 798 64128 134914 65208
rect 880 63848 134914 64128
rect 798 62088 134914 63848
rect 798 61808 134834 62088
rect 798 60728 134914 61808
rect 880 60448 134914 60728
rect 798 58688 134914 60448
rect 798 58408 134834 58688
rect 798 57328 134914 58408
rect 880 57048 134914 57328
rect 798 55288 134914 57048
rect 798 55008 134834 55288
rect 798 53928 134914 55008
rect 880 53648 134914 53928
rect 798 51888 134914 53648
rect 798 51608 134834 51888
rect 798 50528 134914 51608
rect 880 50248 134914 50528
rect 798 48488 134914 50248
rect 798 48208 134834 48488
rect 798 47128 134914 48208
rect 880 46848 134914 47128
rect 798 45088 134914 46848
rect 798 44808 134834 45088
rect 798 43728 134914 44808
rect 880 43448 134914 43728
rect 798 41688 134914 43448
rect 798 41408 134834 41688
rect 798 40328 134914 41408
rect 880 40048 134914 40328
rect 798 38288 134914 40048
rect 798 38008 134834 38288
rect 798 36928 134914 38008
rect 880 36648 134914 36928
rect 798 34888 134914 36648
rect 798 34608 134834 34888
rect 798 33528 134914 34608
rect 880 33248 134914 33528
rect 798 31488 134914 33248
rect 798 31208 134834 31488
rect 798 30128 134914 31208
rect 880 29848 134914 30128
rect 798 28088 134914 29848
rect 798 27808 134834 28088
rect 798 26728 134914 27808
rect 880 26448 134914 26728
rect 798 24688 134914 26448
rect 798 24408 134834 24688
rect 798 23328 134914 24408
rect 880 23048 134914 23328
rect 798 21288 134914 23048
rect 798 21008 134834 21288
rect 798 19928 134914 21008
rect 880 19648 134914 19928
rect 798 17888 134914 19648
rect 798 17608 134834 17888
rect 798 16528 134914 17608
rect 880 16248 134914 16528
rect 798 15168 134914 16248
rect 798 14888 134834 15168
rect 798 13128 134914 14888
rect 880 12848 134914 13128
rect 798 11768 134914 12848
rect 798 11488 134834 11768
rect 798 9728 134914 11488
rect 880 9448 134914 9728
rect 798 8368 134914 9448
rect 798 8088 134834 8368
rect 798 6328 134914 8088
rect 880 6048 134914 6328
rect 798 4968 134914 6048
rect 798 4688 134834 4968
rect 798 2928 134914 4688
rect 880 2648 134914 2928
rect 798 1568 134914 2648
rect 798 1395 134834 1568
<< metal4 >>
rect 4208 2128 4528 135504
rect 4868 2128 5188 135504
rect 34928 2128 35248 135504
rect 35588 2128 35908 135504
rect 65648 2128 65968 135504
rect 66308 2128 66628 135504
rect 96368 2128 96688 135504
rect 97028 2128 97348 135504
rect 127088 2128 127408 135504
rect 127748 2128 128068 135504
<< obsm4 >>
rect 3371 2347 4128 135149
rect 4608 2347 4788 135149
rect 5268 2347 34848 135149
rect 35328 2347 35508 135149
rect 35988 2347 65568 135149
rect 66048 2347 66228 135149
rect 66708 2347 96288 135149
rect 96768 2347 96948 135149
rect 97428 2347 127008 135149
rect 127488 2347 127668 135149
rect 128148 2347 128557 135149
<< metal5 >>
rect 1056 128550 134644 128870
rect 1056 127890 134644 128210
rect 1056 97914 134644 98234
rect 1056 97254 134644 97574
rect 1056 67278 134644 67598
rect 1056 66618 134644 66938
rect 1056 36642 134644 36962
rect 1056 35982 134644 36302
rect 1056 6006 134644 6326
rect 1056 5346 134644 5666
<< labels >>
rlabel metal4 s 4868 2128 5188 135504 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 135504 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 66308 2128 66628 135504 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 97028 2128 97348 135504 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127748 2128 128068 135504 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 134644 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 134644 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 67278 134644 67598 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 97914 134644 98234 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 128550 134644 128870 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 135504 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 135504 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 135504 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 135504 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 135504 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 134644 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 134644 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 66618 134644 66938 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 97254 134644 97574 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 127890 134644 128210 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 110848 800 110968 6 clk
port 3 nsew signal input
rlabel metal3 s 134914 34688 135714 34808 6 input_tdata[0]
port 4 nsew signal input
rlabel metal3 s 134914 21088 135714 21208 6 input_tdata[10]
port 5 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 input_tdata[11]
port 6 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 input_tdata[12]
port 7 nsew signal input
rlabel metal3 s 134914 125808 135714 125928 6 input_tdata[13]
port 8 nsew signal input
rlabel metal3 s 134914 108808 135714 108928 6 input_tdata[14]
port 9 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 input_tdata[15]
port 10 nsew signal input
rlabel metal2 s 104990 137058 105046 137858 6 input_tdata[16]
port 11 nsew signal input
rlabel metal2 s 76654 137058 76710 137858 6 input_tdata[17]
port 12 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 input_tdata[18]
port 13 nsew signal input
rlabel metal3 s 134914 14968 135714 15088 6 input_tdata[19]
port 14 nsew signal input
rlabel metal2 s 117870 137058 117926 137858 6 input_tdata[1]
port 15 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 input_tdata[20]
port 16 nsew signal input
rlabel metal3 s 134914 112208 135714 112328 6 input_tdata[21]
port 17 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 input_tdata[22]
port 18 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 input_tdata[23]
port 19 nsew signal input
rlabel metal2 s 19338 137058 19394 137858 6 input_tdata[24]
port 20 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 input_tdata[25]
port 21 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 input_tdata[26]
port 22 nsew signal input
rlabel metal2 s 70214 137058 70270 137858 6 input_tdata[27]
port 23 nsew signal input
rlabel metal2 s 38014 137058 38070 137858 6 input_tdata[28]
port 24 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 input_tdata[29]
port 25 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 input_tdata[2]
port 26 nsew signal input
rlabel metal3 s 134914 8168 135714 8288 6 input_tdata[30]
port 27 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 input_tdata[31]
port 28 nsew signal input
rlabel metal2 s 89534 137058 89590 137858 6 input_tdata[3]
port 29 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 input_tdata[4]
port 30 nsew signal input
rlabel metal3 s 134914 68688 135714 68808 6 input_tdata[5]
port 31 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 input_tdata[6]
port 32 nsew signal input
rlabel metal3 s 134914 78888 135714 79008 6 input_tdata[7]
port 33 nsew signal input
rlabel metal2 s 57334 137058 57390 137858 6 input_tdata[8]
port 34 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 input_tdata[9]
port 35 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 input_tready
port 36 nsew signal output
rlabel metal2 s 124310 137058 124366 137858 6 input_tvalid
port 37 nsew signal input
rlabel metal2 s 60554 137058 60610 137858 6 load_weight
port 38 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 output_tdata[0]
port 39 nsew signal output
rlabel metal2 s 41234 137058 41290 137858 6 output_tdata[100]
port 40 nsew signal output
rlabel metal3 s 0 124448 800 124568 6 output_tdata[101]
port 41 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 output_tdata[102]
port 42 nsew signal output
rlabel metal2 s 34794 137058 34850 137858 6 output_tdata[103]
port 43 nsew signal output
rlabel metal3 s 134914 61888 135714 62008 6 output_tdata[104]
port 44 nsew signal output
rlabel metal2 s 44454 137058 44510 137858 6 output_tdata[105]
port 45 nsew signal output
rlabel metal3 s 134914 105408 135714 105528 6 output_tdata[106]
port 46 nsew signal output
rlabel metal3 s 134914 85688 135714 85808 6 output_tdata[107]
port 47 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 output_tdata[108]
port 48 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 output_tdata[109]
port 49 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 output_tdata[10]
port 50 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 output_tdata[110]
port 51 nsew signal output
rlabel metal3 s 134914 17688 135714 17808 6 output_tdata[111]
port 52 nsew signal output
rlabel metal3 s 0 134648 800 134768 6 output_tdata[112]
port 53 nsew signal output
rlabel metal3 s 0 83648 800 83768 6 output_tdata[113]
port 54 nsew signal output
rlabel metal2 s 127530 137058 127586 137858 6 output_tdata[114]
port 55 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 output_tdata[115]
port 56 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 output_tdata[116]
port 57 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 output_tdata[117]
port 58 nsew signal output
rlabel metal2 s 130750 137058 130806 137858 6 output_tdata[118]
port 59 nsew signal output
rlabel metal2 s 133970 137058 134026 137858 6 output_tdata[119]
port 60 nsew signal output
rlabel metal2 s 12898 137058 12954 137858 6 output_tdata[11]
port 61 nsew signal output
rlabel metal2 s 63774 137058 63830 137858 6 output_tdata[120]
port 62 nsew signal output
rlabel metal2 s 16118 137058 16174 137858 6 output_tdata[121]
port 63 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 output_tdata[122]
port 64 nsew signal output
rlabel metal3 s 134914 55088 135714 55208 6 output_tdata[123]
port 65 nsew signal output
rlabel metal2 s 86314 137058 86370 137858 6 output_tdata[124]
port 66 nsew signal output
rlabel metal2 s 3238 137058 3294 137858 6 output_tdata[125]
port 67 nsew signal output
rlabel metal2 s 92754 137058 92810 137858 6 output_tdata[126]
port 68 nsew signal output
rlabel metal3 s 134914 72088 135714 72208 6 output_tdata[127]
port 69 nsew signal output
rlabel metal3 s 134914 132608 135714 132728 6 output_tdata[12]
port 70 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 output_tdata[13]
port 71 nsew signal output
rlabel metal2 s 121090 137058 121146 137858 6 output_tdata[14]
port 72 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 output_tdata[15]
port 73 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 output_tdata[16]
port 74 nsew signal output
rlabel metal3 s 0 131248 800 131368 6 output_tdata[17]
port 75 nsew signal output
rlabel metal3 s 134914 122408 135714 122528 6 output_tdata[18]
port 76 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 output_tdata[19]
port 77 nsew signal output
rlabel metal3 s 134914 48288 135714 48408 6 output_tdata[1]
port 78 nsew signal output
rlabel metal2 s 54114 137058 54170 137858 6 output_tdata[20]
port 79 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 output_tdata[21]
port 80 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 output_tdata[22]
port 81 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 output_tdata[23]
port 82 nsew signal output
rlabel metal3 s 134914 102008 135714 102128 6 output_tdata[24]
port 83 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 output_tdata[25]
port 84 nsew signal output
rlabel metal3 s 0 127848 800 127968 6 output_tdata[26]
port 85 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 output_tdata[27]
port 86 nsew signal output
rlabel metal2 s 133970 0 134026 800 6 output_tdata[28]
port 87 nsew signal output
rlabel metal3 s 134914 31288 135714 31408 6 output_tdata[29]
port 88 nsew signal output
rlabel metal2 s 28354 137058 28410 137858 6 output_tdata[2]
port 89 nsew signal output
rlabel metal3 s 134914 58488 135714 58608 6 output_tdata[30]
port 90 nsew signal output
rlabel metal2 s 124310 0 124366 800 6 output_tdata[31]
port 91 nsew signal output
rlabel metal2 s 31574 137058 31630 137858 6 output_tdata[32]
port 92 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 output_tdata[33]
port 93 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 output_tdata[34]
port 94 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 output_tdata[35]
port 95 nsew signal output
rlabel metal2 s 79874 137058 79930 137858 6 output_tdata[36]
port 96 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 output_tdata[37]
port 97 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 output_tdata[38]
port 98 nsew signal output
rlabel metal3 s 134914 119008 135714 119128 6 output_tdata[39]
port 99 nsew signal output
rlabel metal3 s 134914 41488 135714 41608 6 output_tdata[3]
port 100 nsew signal output
rlabel metal2 s 83094 137058 83150 137858 6 output_tdata[40]
port 101 nsew signal output
rlabel metal2 s 101770 137058 101826 137858 6 output_tdata[41]
port 102 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 output_tdata[42]
port 103 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 output_tdata[43]
port 104 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 output_tdata[44]
port 105 nsew signal output
rlabel metal3 s 134914 11568 135714 11688 6 output_tdata[45]
port 106 nsew signal output
rlabel metal2 s 6458 137058 6514 137858 6 output_tdata[46]
port 107 nsew signal output
rlabel metal3 s 134914 98608 135714 98728 6 output_tdata[47]
port 108 nsew signal output
rlabel metal2 s 47674 137058 47730 137858 6 output_tdata[48]
port 109 nsew signal output
rlabel metal2 s 108210 137058 108266 137858 6 output_tdata[49]
port 110 nsew signal output
rlabel metal2 s 9678 137058 9734 137858 6 output_tdata[4]
port 111 nsew signal output
rlabel metal3 s 134914 27888 135714 28008 6 output_tdata[50]
port 112 nsew signal output
rlabel metal3 s 134914 75488 135714 75608 6 output_tdata[51]
port 113 nsew signal output
rlabel metal2 s 50894 137058 50950 137858 6 output_tdata[52]
port 114 nsew signal output
rlabel metal3 s 134914 51688 135714 51808 6 output_tdata[53]
port 115 nsew signal output
rlabel metal3 s 134914 1368 135714 1488 6 output_tdata[54]
port 116 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 output_tdata[55]
port 117 nsew signal output
rlabel metal3 s 134914 95888 135714 96008 6 output_tdata[56]
port 118 nsew signal output
rlabel metal2 s 111430 137058 111486 137858 6 output_tdata[57]
port 119 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 output_tdata[58]
port 120 nsew signal output
rlabel metal3 s 134914 38088 135714 38208 6 output_tdata[59]
port 121 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 output_tdata[5]
port 122 nsew signal output
rlabel metal3 s 134914 4768 135714 4888 6 output_tdata[60]
port 123 nsew signal output
rlabel metal2 s 25134 137058 25190 137858 6 output_tdata[61]
port 124 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 output_tdata[62]
port 125 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 output_tdata[63]
port 126 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 output_tdata[64]
port 127 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 output_tdata[65]
port 128 nsew signal output
rlabel metal3 s 134914 115608 135714 115728 6 output_tdata[66]
port 129 nsew signal output
rlabel metal3 s 134914 82288 135714 82408 6 output_tdata[67]
port 130 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 output_tdata[68]
port 131 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 output_tdata[69]
port 132 nsew signal output
rlabel metal3 s 134914 44888 135714 45008 6 output_tdata[6]
port 133 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 output_tdata[70]
port 134 nsew signal output
rlabel metal3 s 134914 89088 135714 89208 6 output_tdata[71]
port 135 nsew signal output
rlabel metal3 s 134914 129208 135714 129328 6 output_tdata[72]
port 136 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 output_tdata[73]
port 137 nsew signal output
rlabel metal3 s 134914 136008 135714 136128 6 output_tdata[74]
port 138 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 output_tdata[75]
port 139 nsew signal output
rlabel metal3 s 0 104048 800 104168 6 output_tdata[76]
port 140 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 output_tdata[77]
port 141 nsew signal output
rlabel metal2 s 18 0 74 800 6 output_tdata[78]
port 142 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 output_tdata[79]
port 143 nsew signal output
rlabel metal3 s 0 114248 800 114368 6 output_tdata[7]
port 144 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 output_tdata[80]
port 145 nsew signal output
rlabel metal2 s 73434 137058 73490 137858 6 output_tdata[81]
port 146 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 output_tdata[82]
port 147 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 output_tdata[83]
port 148 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 output_tdata[84]
port 149 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 output_tdata[85]
port 150 nsew signal output
rlabel metal2 s 66994 137058 67050 137858 6 output_tdata[86]
port 151 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 output_tdata[87]
port 152 nsew signal output
rlabel metal2 s 114650 137058 114706 137858 6 output_tdata[88]
port 153 nsew signal output
rlabel metal3 s 134914 24488 135714 24608 6 output_tdata[89]
port 154 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 output_tdata[8]
port 155 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 output_tdata[90]
port 156 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 output_tdata[91]
port 157 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 output_tdata[92]
port 158 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 output_tdata[93]
port 159 nsew signal output
rlabel metal3 s 134914 92488 135714 92608 6 output_tdata[94]
port 160 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 output_tdata[95]
port 161 nsew signal output
rlabel metal2 s 98550 137058 98606 137858 6 output_tdata[96]
port 162 nsew signal output
rlabel metal2 s 95974 137058 96030 137858 6 output_tdata[97]
port 163 nsew signal output
rlabel metal2 s 18 137058 74 137858 6 output_tdata[98]
port 164 nsew signal output
rlabel metal2 s 21914 137058 21970 137858 6 output_tdata[99]
port 165 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 output_tdata[9]
port 166 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 output_tready
port 167 nsew signal input
rlabel metal3 s 0 117648 800 117768 6 output_tvalid
port 168 nsew signal output
rlabel metal3 s 134914 65288 135714 65408 6 reset
port 169 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 135714 137858
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 35635690
string GDS_FILE /openlane/designs/tpu/runs/init/results/signoff/top_hardened.magic.gds
string GDS_START 1206826
<< end >>

