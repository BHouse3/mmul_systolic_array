* NGSPICE file created from top_hardened.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s4s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt top_hardened VGND VPWR clk input_tdata[0] input_tdata[10] input_tdata[11]
+ input_tdata[12] input_tdata[13] input_tdata[14] input_tdata[15] input_tdata[16]
+ input_tdata[17] input_tdata[18] input_tdata[19] input_tdata[1] input_tdata[20] input_tdata[21]
+ input_tdata[22] input_tdata[23] input_tdata[24] input_tdata[25] input_tdata[26]
+ input_tdata[27] input_tdata[28] input_tdata[29] input_tdata[2] input_tdata[30] input_tdata[31]
+ input_tdata[3] input_tdata[4] input_tdata[5] input_tdata[6] input_tdata[7] input_tdata[8]
+ input_tdata[9] input_tready input_tvalid load_weight output_tdata[0] output_tdata[100]
+ output_tdata[101] output_tdata[102] output_tdata[103] output_tdata[104] output_tdata[105]
+ output_tdata[106] output_tdata[107] output_tdata[108] output_tdata[109] output_tdata[10]
+ output_tdata[110] output_tdata[111] output_tdata[112] output_tdata[113] output_tdata[114]
+ output_tdata[115] output_tdata[116] output_tdata[117] output_tdata[118] output_tdata[119]
+ output_tdata[11] output_tdata[120] output_tdata[121] output_tdata[122] output_tdata[123]
+ output_tdata[124] output_tdata[125] output_tdata[126] output_tdata[127] output_tdata[12]
+ output_tdata[13] output_tdata[14] output_tdata[15] output_tdata[16] output_tdata[17]
+ output_tdata[18] output_tdata[19] output_tdata[1] output_tdata[20] output_tdata[21]
+ output_tdata[22] output_tdata[23] output_tdata[24] output_tdata[25] output_tdata[26]
+ output_tdata[27] output_tdata[28] output_tdata[29] output_tdata[2] output_tdata[30]
+ output_tdata[31] output_tdata[32] output_tdata[33] output_tdata[34] output_tdata[35]
+ output_tdata[36] output_tdata[37] output_tdata[38] output_tdata[39] output_tdata[3]
+ output_tdata[40] output_tdata[41] output_tdata[42] output_tdata[43] output_tdata[44]
+ output_tdata[45] output_tdata[46] output_tdata[47] output_tdata[48] output_tdata[49]
+ output_tdata[4] output_tdata[50] output_tdata[51] output_tdata[52] output_tdata[53]
+ output_tdata[54] output_tdata[55] output_tdata[56] output_tdata[57] output_tdata[58]
+ output_tdata[59] output_tdata[5] output_tdata[60] output_tdata[61] output_tdata[62]
+ output_tdata[63] output_tdata[64] output_tdata[65] output_tdata[66] output_tdata[67]
+ output_tdata[68] output_tdata[69] output_tdata[6] output_tdata[70] output_tdata[71]
+ output_tdata[72] output_tdata[73] output_tdata[74] output_tdata[75] output_tdata[76]
+ output_tdata[77] output_tdata[78] output_tdata[79] output_tdata[7] output_tdata[80]
+ output_tdata[81] output_tdata[82] output_tdata[83] output_tdata[84] output_tdata[85]
+ output_tdata[86] output_tdata[87] output_tdata[88] output_tdata[89] output_tdata[8]
+ output_tdata[90] output_tdata[91] output_tdata[92] output_tdata[93] output_tdata[94]
+ output_tdata[95] output_tdata[96] output_tdata[97] output_tdata[98] output_tdata[99]
+ output_tdata[9] output_tready output_tvalid reset
XFILLER_0_236_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18869_ _11292_ _11293_ VGND VGND VPWR VPWR _11294_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_234_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20900_ _02669_ _02670_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__or2b_1
XFILLER_0_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21880_ _03453_ _03580_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20831_ _02603_ _02604_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23550_ clknet_leaf_130_clk _00083_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_20762_ _02454_ _02536_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22501_ net654 _05316_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__or2_1
X_23481_ clknet_leaf_136_clk net338 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[71\]
+ sky130_fd_sc_hd__dfxtp_1
X_20693_ _02466_ _02469_ _02471_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__and3_1
XFILLER_0_212_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22432_ _04080_ _04079_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22363_ net711 _05316_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24102_ clknet_leaf_15_clk _00635_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_21314_ top_inst.grid_inst.data_path_wires\[17\]\[0\] _02897_ VGND VGND VPWR VPWR
+ _03052_ sky130_fd_sc_hd__and2b_1
XFILLER_0_131_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22294_ _03979_ _03980_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24033_ clknet_leaf_41_clk _00566_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold340 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[18\] VGND
+ VGND VPWR VPWR net522 sky130_fd_sc_hd__dlygate4sd3_1
X_21245_ _02955_ _02957_ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__or2b_1
Xhold351 top_inst.deskew_buff_inst.col_input\[116\] VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold362 top_inst.deskew_buff_inst.col_input\[79\] VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold373 _00237_ VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[13\] VGND
+ VGND VPWR VPWR net566 sky130_fd_sc_hd__dlygate4sd3_1
X_21176_ _02917_ _02918_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_1111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold395 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[9\] VGND
+ VGND VPWR VPWR net577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20127_ _01934_ _01938_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__xor2_2
XFILLER_0_102_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_217_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20058_ _01562_ _01872_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__nor2_1
XFILLER_0_198_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11900_ net652 _04956_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__or2_1
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ _05653_ _05658_ _05651_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__o21a_1
XFILLER_0_169_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23817_ clknet_leaf_73_clk _00350_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11831_ net599 _04917_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__or2_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _07242_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ net666 _04860_ _04879_ _04875_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__o211a_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23748_ clknet_leaf_122_clk _00281_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13501_ top_inst.grid_inst.data_path_wires\[2\]\[1\] top_inst.grid_inst.data_path_wires\[2\]\[0\]
+ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _06252_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[5\] _07060_ _07173_
+ _07174_ VGND VGND VPWR VPWR _07175_ sky130_fd_sc_hd__and4_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23679_ clknet_leaf_116_clk net597 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16220_ _08802_ _08803_ VGND VGND VPWR VPWR _08804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13432_ _06196_ _05262_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_920 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16151_ _08722_ _08736_ _08737_ VGND VGND VPWR VPWR _08738_ sky130_fd_sc_hd__nand3_2
XFILLER_0_84_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13363_ _06133_ _06135_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer7 _11681_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_148_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15102_ _07750_ _07751_ VGND VGND VPWR VPWR _07752_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12314_ net535 _05183_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__or2_1
X_16082_ _08152_ _08663_ _08680_ _08666_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__o211a_1
X_13294_ _06068_ _06069_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__nor2_1
XFILLER_0_210_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19910_ _01718_ _01731_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__xnor2_2
X_15033_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[3\] _05326_ VGND
+ VGND VPWR VPWR _07686_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12245_ _05127_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__buf_2
XFILLER_0_121_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19841_ _01611_ _01663_ _01664_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__and3_1
X_12176_ _05009_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__buf_2
XFILLER_0_236_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19772_ _01566_ _01568_ _01598_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__a21o_1
X_16984_ _08831_ _09538_ VGND VGND VPWR VPWR _09539_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18723_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _11158_ sky130_fd_sc_hd__clkbuf_4
X_15935_ _08543_ _08545_ VGND VGND VPWR VPWR _08546_ sky130_fd_sc_hd__and2_1
XTAP_5160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18654_ _11109_ _11111_ VGND VGND VPWR VPWR _11112_ sky130_fd_sc_hd__xor2_1
XFILLER_0_189_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15866_ _08458_ _08460_ VGND VGND VPWR VPWR _08478_ sky130_fd_sc_hd__nor2_1
XTAP_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14817_ _07415_ _07501_ VGND VGND VPWR VPWR _07503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17605_ _10113_ _10117_ VGND VGND VPWR VPWR _10118_ sky130_fd_sc_hd__xor2_2
XFILLER_0_231_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1042 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18585_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[14\] _10923_ VGND
+ VGND VPWR VPWR _11045_ sky130_fd_sc_hd__and2_1
XFILLER_0_235_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15797_ _08404_ _08410_ VGND VGND VPWR VPWR _08411_ sky130_fd_sc_hd__xor2_1
XFILLER_0_171_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17536_ _10035_ _10046_ _10055_ _10049_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14748_ _07434_ _07435_ VGND VGND VPWR VPWR _07436_ sky130_fd_sc_hd__xor2_1
XFILLER_0_175_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17467_ _09972_ _10002_ VGND VGND VPWR VPWR _10003_ sky130_fd_sc_hd__xnor2_1
X_14679_ _07366_ _07367_ VGND VGND VPWR VPWR _07368_ sky130_fd_sc_hd__and2b_1
XFILLER_0_188_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19206_ _11479_ _11601_ VGND VGND VPWR VPWR _11622_ sky130_fd_sc_hd__nor2_1
X_16418_ _08831_ _08997_ VGND VGND VPWR VPWR _08998_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17398_ _09915_ _09936_ VGND VGND VPWR VPWR _09937_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_172_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19137_ _11553_ _11554_ VGND VGND VPWR VPWR _11555_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16349_ _08929_ VGND VGND VPWR VPWR _08930_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_923 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19068_ _11479_ _11487_ VGND VGND VPWR VPWR _11488_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18019_ _10511_ _10514_ VGND VGND VPWR VPWR _10521_ sky130_fd_sc_hd__or2_1
XFILLER_0_199_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21030_ _02784_ _02794_ _02795_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__nand3_1
XFILLER_0_22_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_1199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_236_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22981_ net602 _04570_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__or2_1
XFILLER_0_242_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21932_ _03641_ _03648_ _06178_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21863_ _03581_ _03582_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23602_ clknet_leaf_104_clk _00135_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20814_ _02562_ _02588_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24582_ clknet_leaf_142_clk _01115_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dfxtp_1
X_21794_ _03516_ _03511_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23533_ clknet_leaf_140_clk net683 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_20745_ _02465_ _02520_ _02521_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__and3_1
XFILLER_0_212_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23464_ net608 _04859_ _04854_ _06180_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__o211a_1
X_20676_ _02419_ _02451_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22415_ _04097_ _04098_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__or2_1
X_23395_ net729 _04655_ _04817_ _04808_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22346_ _03709_ _03690_ _03990_ _04031_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22277_ _03913_ _03911_ VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__and2b_1
XFILLER_0_103_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12030_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[17\] _05023_
+ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__or2_1
X_24016_ clknet_leaf_52_clk _00549_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_21228_ top_inst.grid_inst.data_path_wires\[17\]\[1\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[17\]\[2\]
+ VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold170 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[22\] VGND
+ VGND VPWR VPWR net352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _00012_ VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold192 _00176_ VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21159_ _02864_ _02862_ _02885_ _02883_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__nand4_2
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13981_ _06698_ _06699_ VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_244_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15720_ _08284_ _08291_ VGND VGND VPWR VPWR _08336_ sky130_fd_sc_hd__or2b_1
X_12932_ _04865_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_198_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _08268_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12863_ _05632_ _05669_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__nor2_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[7\] _07292_ _07069_
+ _07087_ VGND VGND VPWR VPWR _07293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11814_ net933 _04898_ _04908_ _04902_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ _10818_ _10821_ VGND VGND VPWR VPWR _10835_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _08199_ _08201_ VGND VGND VPWR VPWR _08202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12794_ _05569_ _05570_ _05568_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__o21a_1
XFILLER_0_185_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _05399_ _09863_ VGND VGND VPWR VPWR _09864_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14533_ _07117_ _07225_ VGND VGND VPWR VPWR _07226_ sky130_fd_sc_hd__and2_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11745_ net36 VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__buf_8
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17252_ _09791_ _09797_ VGND VGND VPWR VPWR _09798_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14464_ _07156_ _07157_ _07057_ VGND VGND VPWR VPWR _07159_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16203_ _08762_ _08786_ _08265_ VGND VGND VPWR VPWR _08788_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13415_ _06184_ _05262_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__or2_1
X_17183_ _09729_ _09730_ _09623_ VGND VGND VPWR VPWR _09732_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_180_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14395_ _07062_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[0\] _07061_
+ VGND VGND VPWR VPWR _07094_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16134_ _06848_ _08720_ _08721_ _08692_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__o211a_1
X_13346_ _06084_ _06088_ _06119_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16065_ _08139_ _08663_ _08668_ _08666_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__o211a_1
X_13277_ _06016_ _06051_ _05980_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15016_ _07606_ _07633_ _07631_ _07608_ VGND VGND VPWR VPWR _07669_ sky130_fd_sc_hd__a22o_1
X_12228_ net812 _05137_ _05145_ _05141_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19824_ _01556_ _01591_ _01648_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__or3b_4
XFILLER_0_236_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12159_ net775 _05097_ _05105_ _05101_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19755_ _01580_ _01581_ _01569_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__a21o_1
XFILLER_0_237_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_208_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16967_ _09518_ _09519_ _09520_ VGND VGND VPWR VPWR _09522_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18706_ _10592_ _11142_ _11146_ _11137_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__o211a_1
X_15918_ _08516_ _08492_ _08527_ VGND VGND VPWR VPWR _08529_ sky130_fd_sc_hd__nand3_1
X_16898_ _09410_ _09446_ VGND VGND VPWR VPWR _09454_ sky130_fd_sc_hd__or2b_1
X_19686_ _01428_ _01467_ _01468_ _01511_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__or4b_4
XFILLER_0_91_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15849_ _08415_ _08419_ _08417_ VGND VGND VPWR VPWR _08462_ sky130_fd_sc_hd__a21oi_1
X_18637_ net1067 _10616_ _11095_ _10620_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__o211a_1
XFILLER_0_232_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18568_ _10974_ _10989_ _11028_ VGND VGND VPWR VPWR _11029_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17519_ _10022_ _08681_ _10043_ _10024_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18499_ _10946_ _10947_ VGND VGND VPWR VPWR _10961_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20530_ _02274_ _02281_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20461_ _02193_ _02194_ _02244_ _02245_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__a211o_1
XFILLER_0_172_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22200_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[7\] _03852_ _03853_
+ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__a21boi_2
X_23180_ net723 _04685_ _04696_ _04691_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20392_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _02178_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22131_ _03709_ _03682_ top_inst.grid_inst.data_path_wires\[18\]\[0\] _03711_ VGND
+ VGND VPWR VPWR _03822_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_140_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22062_ _05312_ _03753_ _03754_ _03755_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__a31o_1
XTAP_6619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_220_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21013_ _05405_ _02779_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__nor2_1
XTAP_5907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22964_ net602 _04562_ _04571_ _04564_ VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__o211a_1
XFILLER_0_241_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21915_ _03576_ _03630_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22895_ top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[4\] _04530_ VGND
+ VGND VPWR VPWR _04532_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24634_ clknet_leaf_26_clk _01167_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[110\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21846_ _03539_ _03565_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__or2_1
XFILLER_0_194_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24565_ clknet_leaf_137_clk _01098_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_194_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21777_ _03499_ _03500_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23516_ clknet_leaf_138_clk _00049_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20728_ _02495_ _02505_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24496_ clknet_leaf_126_clk _01029_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_135_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23447_ net460 _04835_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20659_ _02188_ _02438_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__and2b_1
XFILLER_0_190_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_1306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13200_ _05750_ top_inst.grid_inst.data_path_wires\[1\]\[5\] _05765_ _05763_ VGND
+ VGND VPWR VPWR _05978_ sky130_fd_sc_hd__and4_1
XFILLER_0_151_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14180_ _06891_ _06892_ VGND VGND VPWR VPWR _06893_ sky130_fd_sc_hd__nor2_1
X_23378_ net52 _04805_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13131_ _05901_ _05910_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22329_ _03978_ _03981_ _04014_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_143_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13062_ _05818_ _05843_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__or2_1
XFILLER_0_237_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12013_ net883 _05018_ _05021_ _05022_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__o211a_1
X_17870_ _10335_ _10375_ VGND VGND VPWR VPWR _10376_ sky130_fd_sc_hd__nor2_2
XFILLER_0_40_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16821_ _09361_ _09186_ _09191_ _09213_ VGND VGND VPWR VPWR _09379_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_191_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16752_ _09302_ _09303_ _09310_ VGND VGND VPWR VPWR _09312_ sky130_fd_sc_hd__a21oi_1
X_19540_ _01312_ _01320_ _01319_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__a21bo_1
X_13964_ _05260_ VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15703_ _08147_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[2\] _08317_
+ _08318_ VGND VGND VPWR VPWR _08319_ sky130_fd_sc_hd__a22o_1
X_12915_ _05718_ _05406_ _05719_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__or3b_1
XFILLER_0_214_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16683_ _08831_ _09245_ VGND VGND VPWR VPWR _09246_ sky130_fd_sc_hd__and2_1
X_19471_ _01300_ _01304_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_232_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13895_ _06190_ _06192_ _06629_ _06446_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15634_ _08250_ _08251_ VGND VGND VPWR VPWR _08252_ sky130_fd_sc_hd__nand2_1
X_18422_ _10595_ _10602_ _10849_ _10850_ VGND VGND VPWR VPWR _10886_ sky130_fd_sc_hd__a31o_1
X_12846_ _05651_ _05652_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _10775_ _10752_ VGND VGND VPWR VPWR _10819_ sky130_fd_sc_hd__or2b_1
XFILLER_0_111_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15565_ _08184_ _08185_ VGND VGND VPWR VPWR _08186_ sky130_fd_sc_hd__nand2_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _05579_ _05580_ _05584_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17304_ _09830_ _09831_ _09847_ VGND VGND VPWR VPWR _09848_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_173_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14516_ _07175_ _07207_ _07208_ VGND VGND VPWR VPWR _07209_ sky130_fd_sc_hd__nand3_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_230_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18284_ _10717_ _10721_ _10750_ VGND VGND VPWR VPWR _10751_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_232_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15496_ top_inst.grid_inst.data_path_wires\[7\]\[0\] VGND VGND VPWR VPWR _08135_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17235_ _09761_ _09781_ VGND VGND VPWR VPWR _09782_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14447_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[3\] _07119_ _07120_
+ VGND VGND VPWR VPWR _07142_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_226_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17166_ _09697_ _09715_ VGND VGND VPWR VPWR _09716_ sky130_fd_sc_hd__and2_1
XFILLER_0_142_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_226_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14378_ _05290_ _07078_ _07080_ _06684_ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_243_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold906 top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[15\] VGND VGND
+ VPWR VPWR net1088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold917 top_inst.deskew_buff_inst.col_input\[25\] VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__dlygate4sd3_1
X_16117_ _08703_ _08704_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[1\]
+ VGND VGND VPWR VPWR _08706_ sky130_fd_sc_hd__a21o_1
Xhold928 top_inst.axis_in_inst.inbuf_bus\[23\] VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ _06065_ _06103_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__xnor2_1
X_17097_ _09594_ _09608_ _09607_ VGND VGND VPWR VPWR _09649_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16048_ _08640_ _08654_ VGND VGND VPWR VPWR _08655_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19807_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[14\] _01395_ _01396_
+ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17999_ _10498_ _10501_ VGND VGND VPWR VPWR _10502_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19738_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[12\] _01395_ _01396_
+ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__a21o_1
XFILLER_0_237_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19669_ _01444_ _01452_ _01451_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_133_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21700_ _03425_ _03426_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22680_ _04352_ _04353_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__nor2_1
XFILLER_0_177_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_946 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21631_ _03359_ _03360_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__and2b_1
XFILLER_0_158_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24350_ clknet_leaf_24_clk _00883_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[109\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21562_ _03290_ _03293_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__xor2_2
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23301_ net687 _04752_ _04764_ _04756_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20513_ _02294_ _02295_ _02296_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__nand3_2
XFILLER_0_160_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21493_ _03200_ _03226_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__xor2_2
X_24281_ clknet_leaf_11_clk _00814_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23232_ net699 _04713_ _04725_ _04717_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__o211a_1
X_20444_ _02178_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_244_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_209_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23163_ _04657_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20375_ _02143_ _02160_ _02161_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__nor3_2
XFILLER_0_101_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22114_ _03805_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__clkbuf_1
X_23094_ _09787_ _04645_ _04867_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__a21oi_1
XTAP_6405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22045_ _03703_ _03682_ _03680_ _03705_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__a22o_1
XTAP_6449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23996_ clknet_4_14__leaf_clk _00529_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1034 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22947_ net662 _04548_ _04561_ _04551_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12700_ _05509_ _05510_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13680_ _06371_ _06424_ _06425_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_57_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22878_ _10583_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_151_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12631_ _05423_ _05426_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__and2_1
X_24617_ clknet_leaf_32_clk _01150_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_151_1376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21829_ _03536_ _03529_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__and2b_1
XFILLER_0_13_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15350_ _07992_ _07993_ VGND VGND VPWR VPWR _07994_ sky130_fd_sc_hd__or2_1
X_12562_ _05362_ _05365_ _05367_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__or3_1
XFILLER_0_183_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24548_ clknet_leaf_100_clk _01081_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_53_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14301_ _06981_ _07010_ VGND VGND VPWR VPWR _07011_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15281_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[10\] _07845_ VGND
+ VGND VPWR VPWR _07927_ sky130_fd_sc_hd__xnor2_2
X_24479_ clknet_leaf_55_clk _01012_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12493_ _05311_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__buf_8
XFILLER_0_227_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17020_ _09499_ _09526_ _09525_ VGND VGND VPWR VPWR _09574_ sky130_fd_sc_hd__a21bo_1
X_14232_ _06632_ _06898_ _06899_ _06860_ VGND VGND VPWR VPWR _06944_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_135_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14163_ _06830_ _06876_ _06827_ VGND VGND VPWR VPWR _06877_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13114_ _05855_ _05893_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__xor2_1
X_14094_ _06807_ _06808_ VGND VGND VPWR VPWR _06809_ sky130_fd_sc_hd__nor2_1
X_18971_ _11388_ _11392_ VGND VGND VPWR VPWR _11393_ sky130_fd_sc_hd__xor2_1
XFILLER_0_238_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ top_inst.grid_inst.data_path_wires\[1\]\[3\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[2\]
+ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__and2_1
X_17922_ _10425_ _10426_ VGND VGND VPWR VPWR _10427_ sky130_fd_sc_hd__xnor2_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_2__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_4_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17853_ _10324_ _10359_ VGND VGND VPWR VPWR _10360_ sky130_fd_sc_hd__nand2_1
X_16804_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[6\] _09325_ _09326_
+ VGND VGND VPWR VPWR _09362_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_156_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14996_ _07648_ _07649_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[1\]
+ VGND VGND VPWR VPWR _07651_ sky130_fd_sc_hd__a21o_1
X_17784_ top_inst.grid_inst.data_path_wires\[11\]\[5\] _10052_ _10050_ _10037_ VGND
+ VGND VPWR VPWR _10292_ sky130_fd_sc_hd__a22o_1
XFILLER_0_234_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19523_ _01351_ _01355_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16735_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[4\] _09274_ _09275_
+ VGND VGND VPWR VPWR _09295_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_163_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13947_ _06666_ _06667_ _05328_ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16666_ _09228_ _09229_ _08181_ VGND VGND VPWR VPWR _09230_ sky130_fd_sc_hd__o21ai_1
X_19454_ _01221_ _01259_ _01287_ _01288_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13878_ net1074 _06169_ _06616_ _06617_ _06180_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__o221a_1
XFILLER_0_88_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18405_ _10867_ _10869_ VGND VGND VPWR VPWR _10870_ sky130_fd_sc_hd__xnor2_1
X_15617_ _08233_ _08234_ _07057_ VGND VGND VPWR VPWR _08236_ sky130_fd_sc_hd__a21o_1
X_12829_ _05619_ _05620_ _05622_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__or3b_1
XFILLER_0_201_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16597_ _09149_ _09171_ _04870_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19385_ _01218_ _01219_ _01220_ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_243_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18336_ _10585_ _10610_ VGND VGND VPWR VPWR _10802_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15548_ _08152_ _07639_ _08171_ _08166_ VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__o211a_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18267_ _10723_ _10734_ VGND VGND VPWR VPWR _10735_ sky130_fd_sc_hd__nand2_1
X_15479_ _08116_ _08118_ VGND VGND VPWR VPWR _08120_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17218_ _09741_ _09744_ _09764_ _07439_ VGND VGND VPWR VPWR _09766_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18198_ _10646_ _10667_ VGND VGND VPWR VPWR _10668_ sky130_fd_sc_hd__xor2_2
XFILLER_0_170_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold703 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[17\] VGND
+ VGND VPWR VPWR net885 sky130_fd_sc_hd__dlygate4sd3_1
X_17149_ _09681_ _09682_ VGND VGND VPWR VPWR _09699_ sky130_fd_sc_hd__or2_1
Xhold714 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[6\] VGND
+ VGND VPWR VPWR net896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold725 top_inst.deskew_buff_inst.col_input\[19\] VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 top_inst.axis_in_inst.inbuf_bus\[19\] VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold747 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[31\] VGND
+ VGND VPWR VPWR net929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20160_ top_inst.deskew_buff_inst.col_input\[30\] _11723_ _01969_ _01970_ VGND VGND
+ VPWR VPWR _01971_ sky130_fd_sc_hd__a22o_1
Xhold758 top_inst.axis_out_inst.out_buff_data\[68\] VGND VGND VPWR VPWR net940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 top_inst.axis_in_inst.inbuf_bus\[2\] VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20091_ _01903_ _01904_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__nor2_1
XFILLER_0_196_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_224_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23850_ clknet_leaf_68_clk _00383_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22801_ _04388_ _04446_ _04468_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23781_ clknet_leaf_65_clk _00314_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20993_ _02735_ _02757_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__or2b_1
XFILLER_0_211_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22732_ _04377_ _04403_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22663_ _04319_ _04336_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_220_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24402_ clknet_leaf_57_clk net770 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].output_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_21614_ top_inst.deskew_buff_inst.col_input\[78\] _05731_ _03343_ _03344_ VGND VGND
+ VPWR VPWR _03345_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22594_ _04261_ _04270_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_1360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24333_ clknet_leaf_5_clk _00866_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21545_ _03275_ _03272_ _03276_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_209_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_141_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_141_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_173_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24264_ clknet_leaf_105_clk _00797_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21476_ _03135_ _03209_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23215_ _04690_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_1418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20427_ _02210_ _02211_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_181_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24195_ clknet_leaf_15_clk _00728_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23146_ net618 _04671_ _04676_ _04675_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20358_ _01986_ _02020_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[0\]
+ top_inst.grid_inst.data_path_wires\[16\]\[6\] VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23077_ net18 _04628_ _04636_ _04632_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__o211a_1
X_20289_ top_inst.grid_inst.data_path_wires\[16\]\[3\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[1\]
+ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__and2_1
XTAP_6246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22028_ _03722_ _03723_ _05732_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__a21o_1
XFILLER_0_228_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14850_ _07527_ _07502_ _07534_ VGND VGND VPWR VPWR _07535_ sky130_fd_sc_hd__o21ba_1
XTAP_5578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold74 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[27\] VGND
+ VGND VPWR VPWR net256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_242_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold85 _00163_ VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_243_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold96 top_inst.deskew_buff_inst.col_input\[47\] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13801_ _06505_ _06509_ _06503_ VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_230_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14781_ _07456_ _07457_ _07466_ VGND VGND VPWR VPWR _07468_ sky130_fd_sc_hd__nand3_1
XTAP_4888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11993_ net737 _05004_ _05011_ _05008_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__o211a_1
X_23979_ clknet_leaf_87_clk _00512_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_16520_ _09095_ _09096_ VGND VGND VPWR VPWR _09097_ sky130_fd_sc_hd__nor2_1
XFILLER_0_230_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13732_ _06474_ _06476_ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__nor2_1
Xclkbuf_4_10__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_4_10__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_196_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16451_ _08976_ _08979_ _09029_ VGND VGND VPWR VPWR _09030_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13663_ _06408_ VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15402_ _08005_ _08044_ VGND VGND VPWR VPWR _08045_ sky130_fd_sc_hd__nor2_1
X_12614_ _05423_ _05426_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__xor2_1
XFILLER_0_186_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19170_ _11586_ VGND VGND VPWR VPWR _11587_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16382_ _08960_ _08961_ VGND VGND VPWR VPWR _08962_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13594_ top_inst.grid_inst.data_path_wires\[2\]\[6\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[2\]\[7\]
+ VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__a22o_1
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18121_ _10599_ _10046_ _10601_ _10594_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15333_ _07976_ _07977_ VGND VGND VPWR VPWR _07978_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12545_ _05358_ _05359_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_132_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_132_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_124_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18052_ _10546_ _10552_ VGND VGND VPWR VPWR _10553_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15264_ _07615_ _07640_ _07824_ _07613_ VGND VGND VPWR VPWR _07910_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12476_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _05298_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17003_ _09554_ net221 _09556_ VGND VGND VPWR VPWR _09557_ sky130_fd_sc_hd__nand3_1
X_14215_ _06652_ top_inst.grid_inst.data_path_wires\[3\]\[5\] _06925_ VGND VGND VPWR
+ VPWR _06927_ sky130_fd_sc_hd__and3_1
XFILLER_0_151_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_5 _07816_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15195_ top_inst.grid_inst.data_path_wires\[6\]\[7\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _07843_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_870 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_240_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_238_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14146_ _06635_ _06643_ VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__nand2_2
XFILLER_0_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14077_ _06739_ _06748_ VGND VGND VPWR VPWR _06793_ sky130_fd_sc_hd__or2_1
X_18954_ _11328_ _11329_ _11376_ VGND VGND VPWR VPWR _11377_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13028_ top_inst.grid_inst.data_path_wires\[1\]\[1\] top_inst.grid_inst.data_path_wires\[1\]\[0\]
+ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _05811_ sky130_fd_sc_hd__and3_1
X_17905_ _10374_ _10390_ _10409_ VGND VGND VPWR VPWR _10410_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_197_1376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18885_ top_inst.grid_inst.data_path_wires\[13\]\[4\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[3\]
+ _11138_ _11158_ VGND VGND VPWR VPWR _11309_ sky130_fd_sc_hd__a22o_1
XTAP_6780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17836_ _10339_ _10342_ VGND VGND VPWR VPWR _10343_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_238_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer17 _09721_ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer28 _01384_ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__buf_1
X_17767_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[8\] _09496_ _10274_
+ _10275_ VGND VGND VPWR VPWR _10276_ sky130_fd_sc_hd__a22o_1
Xrebuffer39 _09555_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14979_ _07637_ _07075_ VGND VGND VPWR VPWR _07638_ sky130_fd_sc_hd__or2_1
XFILLER_0_234_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19506_ _01338_ _01339_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__or2b_1
X_16718_ _09276_ _09277_ _09255_ VGND VGND VPWR VPWR _09279_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17698_ _10035_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[2\] _10205_
+ _10206_ VGND VGND VPWR VPWR _10208_ sky130_fd_sc_hd__nand4_1
X_19437_ _11688_ _11696_ _01270_ _01271_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__nand4_2
XFILLER_0_130_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16649_ _05269_ _09215_ VGND VGND VPWR VPWR _09216_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19368_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[4\] _01203_ _01204_
+ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18319_ _10641_ _10785_ VGND VGND VPWR VPWR _10786_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_123_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_123_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19299_ _05755_ _11696_ _11698_ _11641_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21330_ _03066_ _03067_ top_inst.deskew_buff_inst.col_input\[71\] _05354_ VGND VGND
+ VPWR VPWR _03068_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_128_1131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold500 top_inst.deskew_buff_inst.col_input\[91\] VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__clkdlybuf4s25_1
X_21261_ top_inst.grid_inst.data_path_wires\[17\]\[5\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[1\]
+ _02882_ top_inst.grid_inst.data_path_wires\[17\]\[6\] VGND VGND VPWR VPWR _03000_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold511 top_inst.axis_out_inst.out_buff_data\[51\] VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[3\] VGND VGND
+ VPWR VPWR net704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[0\] VGND VGND
+ VPWR VPWR net715 sky130_fd_sc_hd__dlygate4sd3_1
X_23000_ top_inst.skew_buff_inst.row\[0\].output_reg\[1\] _04583_ VGND VGND VPWR VPWR
+ _04592_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20212_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _02011_ sky130_fd_sc_hd__clkbuf_4
Xhold544 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[23\] VGND
+ VGND VPWR VPWR net726 sky130_fd_sc_hd__dlygate4sd3_1
X_21192_ _02932_ _02933_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold555 top_inst.deskew_buff_inst.col_input\[32\] VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__buf_1
Xhold566 top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[31\] VGND VGND
+ VPWR VPWR net748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[20\] VGND
+ VGND VPWR VPWR net759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 _00935_ VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__dlygate4sd3_1
X_20143_ _01563_ _01952_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold599 top_inst.axis_out_inst.out_buff_data\[97\] VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20074_ _11722_ _01888_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__and2_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23902_ clknet_leaf_52_clk _00435_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23833_ clknet_leaf_93_clk _00366_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23764_ clknet_leaf_66_clk _00297_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20976_ _02466_ _02742_ _02743_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__and3_1
XFILLER_0_178_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22715_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[25\] _03937_ VGND
+ VGND VPWR VPWR _04387_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23695_ clknet_leaf_119_clk _00228_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22646_ _04296_ _04321_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22577_ _04188_ _04254_ _04255_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_118_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_114_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24316_ clknet_leaf_1_clk _00849_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[91\]
+ sky130_fd_sc_hd__dfxtp_1
X_12330_ net345 _05196_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__or2_1
X_21528_ _03210_ _03260_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24247_ clknet_leaf_108_clk _00780_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_12261_ net925 _05151_ _05163_ _05155_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__o211a_1
X_21459_ _03190_ _03192_ _10831_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__o21a_1
X_14000_ top_inst.grid_inst.data_path_wires\[3\]\[4\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[3\]\[5\]
+ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_142_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24178_ clknet_leaf_29_clk _00711_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12192_ top_inst.axis_out_inst.out_buff_data\[23\] _05115_ VGND VGND VPWR VPWR _05124_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_222_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput42 net42 VGND VGND VPWR VPWR output_tdata[103] sky130_fd_sc_hd__clkbuf_4
XTAP_6010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput53 net53 VGND VGND VPWR VPWR output_tdata[113] sky130_fd_sc_hd__clkbuf_4
X_23129_ net686 _04656_ _04666_ _04662_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__o211a_1
XTAP_6021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput64 net64 VGND VGND VPWR VPWR output_tdata[123] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_235_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput75 net75 VGND VGND VPWR VPWR output_tdata[18] sky130_fd_sc_hd__buf_2
XTAP_6043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput86 net86 VGND VGND VPWR VPWR output_tdata[28] sky130_fd_sc_hd__clkbuf_4
XTAP_6054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput97 net97 VGND VGND VPWR VPWR output_tdata[38] sky130_fd_sc_hd__clkbuf_4
XTAP_6065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15951_ _08559_ _08560_ VGND VGND VPWR VPWR _08561_ sky130_fd_sc_hd__nor2_1
XTAP_6076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14902_ _07582_ _07584_ VGND VGND VPWR VPWR _07585_ sky130_fd_sc_hd__xnor2_1
XTAP_6098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18670_ _11090_ _11112_ VGND VGND VPWR VPWR _11127_ sky130_fd_sc_hd__and2b_1
X_15882_ _08492_ _08493_ VGND VGND VPWR VPWR _08494_ sky130_fd_sc_hd__nand2_1
XTAP_5375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ _10127_ _10132_ VGND VGND VPWR VPWR _10133_ sky130_fd_sc_hd__xnor2_2
X_14833_ _07483_ _07480_ _07517_ _07439_ VGND VGND VPWR VPWR _07519_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_1056 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14764_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[12\] _07281_ VGND
+ VGND VPWR VPWR _07451_ sky130_fd_sc_hd__xnor2_1
XTAP_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ _10066_ _10067_ _10061_ VGND VGND VPWR VPWR _10068_ sky130_fd_sc_hd__a21o_1
XTAP_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ net1101 _04996_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__or2_1
XFILLER_0_230_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16503_ _09045_ _09046_ VGND VGND VPWR VPWR _09080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13715_ _06196_ _06458_ _06459_ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_233_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17483_ _09625_ _09919_ _10016_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[27\]
+ VGND VGND VPWR VPWR _10017_ sky130_fd_sc_hd__a31o_1
XFILLER_0_156_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14695_ _07334_ _07336_ VGND VGND VPWR VPWR _07384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19222_ _11620_ _11637_ VGND VGND VPWR VPWR _11638_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16434_ _08961_ _08963_ _08960_ VGND VGND VPWR VPWR _09013_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_2_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13646_ _06383_ _06392_ VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16365_ _08892_ _08904_ _08945_ VGND VGND VPWR VPWR _08946_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19153_ _11569_ _11570_ VGND VGND VPWR VPWR _11571_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_105_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13577_ _05886_ _06325_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15316_ _07621_ _07637_ VGND VGND VPWR VPWR _07961_ sky130_fd_sc_hd__nand2_1
X_18104_ top_inst.grid_inst.data_path_wires\[12\]\[5\] VGND VGND VPWR VPWR _10589_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12528_ _05341_ _05343_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__xor2_1
X_16296_ _08875_ _08877_ VGND VGND VPWR VPWR _08878_ sky130_fd_sc_hd__nor2_2
X_19084_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[11\] _10364_ _11502_
+ _11503_ _11228_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__o221a_1
XFILLER_0_125_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_240_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15247_ _07839_ _07837_ VGND VGND VPWR VPWR _07894_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18035_ _10534_ _10535_ VGND VGND VPWR VPWR _10537_ sky130_fd_sc_hd__nand2_1
X_12459_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _05284_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_239_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15178_ _07823_ _07825_ VGND VGND VPWR VPWR _07826_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14129_ _06801_ _06802_ _06843_ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_239_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19986_ _01561_ _01802_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18937_ _11313_ _11319_ _11359_ VGND VGND VPWR VPWR _11360_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_1094 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18868_ _11203_ _11224_ _11250_ _11254_ VGND VGND VPWR VPWR _11293_ sky130_fd_sc_hd__o31a_1
XFILLER_0_206_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17819_ _10313_ _10282_ VGND VGND VPWR VPWR _10326_ sky130_fd_sc_hd__or2b_1
XFILLER_0_179_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18799_ _11224_ _11225_ VGND VGND VPWR VPWR _11226_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20830_ _02528_ _02595_ _02602_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__nand3_1
XFILLER_0_72_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20761_ _02385_ _02388_ _02537_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_175_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_523 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22500_ _04160_ _04156_ _04180_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23480_ clknet_leaf_136_clk net361 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20692_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[14\] _02470_ VGND
+ VGND VPWR VPWR _02471_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22431_ _04093_ _04114_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22362_ _04012_ _04008_ _04046_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24101_ clknet_leaf_15_clk _00634_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_103_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21313_ top_inst.grid_inst.data_path_wires\[17\]\[1\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__nand2_1
X_22293_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[10\] _03894_ VGND
+ VGND VPWR VPWR _03980_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_206_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24032_ clknet_leaf_53_clk _00565_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold330 top_inst.axis_out_inst.out_buff_data\[100\] VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21244_ _02981_ _02983_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__xnor2_2
Xhold341 _00025_ VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 _01173_ VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 _00054_ VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold374 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[2\] VGND
+ VGND VPWR VPWR net556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[13\] VGND
+ VGND VPWR VPWR net567 sky130_fd_sc_hd__dlygate4sd3_1
X_21175_ _02910_ _02916_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__nand2_1
XFILLER_0_217_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold396 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[1\] VGND VGND
+ VPWR VPWR net578 sky130_fd_sc_hd__dlygate4sd3_1
X_20126_ _01936_ _01937_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__and2b_1
X_20057_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[26\] _01764_ VGND
+ VGND VPWR VPWR _01872_ sky130_fd_sc_hd__xnor2_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1090 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23816_ clknet_leaf_73_clk _00349_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_11830_ net794 _04912_ _04918_ _04916_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__o211a_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11761_ top_inst.axis_out_inst.out_buff_data\[125\] _04877_ VGND VGND VPWR VPWR _04879_
+ sky130_fd_sc_hd__or2_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23747_ clknet_leaf_122_clk net320 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20959_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[21\] _02559_ _02692_
+ _02690_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13500_ _06186_ _06205_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__nand2_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14480_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[2\] _07073_ _07171_
+ _07172_ VGND VGND VPWR VPWR _07174_ sky130_fd_sc_hd__a22o_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23678_ clknet_leaf_117_clk net827 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13431_ _06195_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_180_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22629_ _09787_ _04304_ _04305_ _03929_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16150_ _08723_ _08717_ _08735_ VGND VGND VPWR VPWR _08737_ sky130_fd_sc_hd__nand3_1
XFILLER_0_180_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13362_ _06133_ _06135_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer8 net189 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__buf_6
X_15101_ _07615_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[2\] _07748_
+ _07749_ VGND VGND VPWR VPWR _07751_ sky130_fd_sc_hd__nand4_2
XFILLER_0_224_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12313_ net841 _05191_ _05193_ _05182_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__o211a_1
X_16081_ _08679_ _08674_ VGND VGND VPWR VPWR _08680_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13293_ _06023_ _06027_ _06021_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_161_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15032_ _07682_ _07683_ _07667_ VGND VGND VPWR VPWR _07685_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12244_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[13\] _05143_
+ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19840_ _01663_ _01664_ _01611_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12175_ net323 _05110_ _05113_ _05114_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19771_ _01562_ _01567_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__nor2_1
X_16983_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[10\] _09496_ _09535_
+ _09537_ VGND VGND VPWR VPWR _09538_ sky130_fd_sc_hd__a22o_1
XFILLER_0_236_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18722_ _11138_ _10607_ _11157_ _11137_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__o211a_1
XTAP_5150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15934_ _08503_ _08504_ _08544_ VGND VGND VPWR VPWR _08545_ sky130_fd_sc_hd__a21bo_1
XTAP_5161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18653_ _11085_ _11086_ _11110_ VGND VGND VPWR VPWR _11111_ sky130_fd_sc_hd__a21oi_1
XTAP_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15865_ _08463_ _08465_ VGND VGND VPWR VPWR _08477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_235_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17604_ _10114_ _10116_ VGND VGND VPWR VPWR _10117_ sky130_fd_sc_hd__xor2_2
XFILLER_0_8_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14816_ _07415_ _07501_ VGND VGND VPWR VPWR _07502_ sky130_fd_sc_hd__and2_1
XFILLER_0_204_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_979 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18584_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[13\] _10923_ _10840_
+ VGND VGND VPWR VPWR _11044_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ _08408_ _08409_ VGND VGND VPWR VPWR _08410_ sky130_fd_sc_hd__xor2_1
XFILLER_0_231_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17535_ _10054_ _09199_ VGND VGND VPWR VPWR _10055_ sky130_fd_sc_hd__or2_1
X_14747_ _07363_ _07393_ _07392_ VGND VGND VPWR VPWR _07435_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_153_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11959_ net693 _04982_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14678_ _07328_ _07331_ _07330_ VGND VGND VPWR VPWR _07367_ sky130_fd_sc_hd__o21ai_1
X_17466_ _09936_ _09956_ _09919_ VGND VGND VPWR VPWR _10002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19205_ _11514_ _11592_ _11594_ VGND VGND VPWR VPWR _11621_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16417_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[10\] _08066_ _08995_
+ _08996_ VGND VGND VPWR VPWR _08997_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13629_ top_inst.grid_inst.data_path_wires\[2\]\[5\] _06190_ _06210_ _06208_ VGND
+ VGND VPWR VPWR _06376_ sky130_fd_sc_hd__nand4_1
XFILLER_0_183_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17397_ _09935_ VGND VGND VPWR VPWR _09936_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19136_ _11514_ _11552_ VGND VGND VPWR VPWR _11554_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16348_ top_inst.grid_inst.data_path_wires\[8\]\[6\] top_inst.grid_inst.data_path_wires\[8\]\[5\]
+ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _08929_ sky130_fd_sc_hd__and4_1
XFILLER_0_229_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16279_ _08860_ _08861_ VGND VGND VPWR VPWR _08862_ sky130_fd_sc_hd__xnor2_1
X_19067_ _11485_ _11486_ VGND VGND VPWR VPWR _11487_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18018_ _10486_ _10516_ _10519_ VGND VGND VPWR VPWR _10520_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_120_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19969_ _01786_ _01787_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__nor2_1
XFILLER_0_238_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22980_ net606 _04575_ _04580_ _04577_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__o211a_1
XFILLER_0_241_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21931_ _03549_ _03643_ _03645_ _03647_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__a211o_1
XFILLER_0_241_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21862_ _03453_ _03560_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__nor2_1
XFILLER_0_214_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23601_ clknet_leaf_103_clk net519 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20813_ _02586_ _02587_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24581_ clknet_leaf_139_clk _01114_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21793_ _03495_ _03515_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23532_ clknet_leaf_139_clk net431 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20744_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[16\] _02467_ VGND
+ VGND VPWR VPWR _02521_ sky130_fd_sc_hd__or2_1
XFILLER_0_175_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23463_ top_inst.axis_out_inst.out_buff_data\[119\] _04864_ VGND VGND VPWR VPWR _04854_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_161_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20675_ _02416_ _02422_ _02450_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22414_ _04094_ _04096_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23394_ net61 _04658_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22345_ _03711_ top_inst.grid_inst.data_path_wires\[18\]\[4\] _03988_ VGND VGND VPWR
+ VPWR _04031_ sky130_fd_sc_hd__and3_1
XFILLER_0_143_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22276_ _03945_ _03963_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24015_ clknet_leaf_48_clk _00548_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_103_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold160 _00185_ VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__dlygate4sd3_1
X_21227_ top_inst.grid_inst.data_path_wires\[17\]\[2\] top_inst.grid_inst.data_path_wires\[17\]\[1\]
+ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[4\] VGND VGND VPWR VPWR
+ _02967_ sky130_fd_sc_hd__and3_1
XFILLER_0_143_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold171 _00189_ VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 top_inst.axis_out_inst.out_buff_data\[66\] VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold193 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[29\] VGND
+ VGND VPWR VPWR net375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21158_ top_inst.grid_inst.data_path_wires\[17\]\[0\] _02885_ _02883_ _02864_ VGND
+ VGND VPWR VPWR _02902_ sky130_fd_sc_hd__a22o_1
XFILLER_0_217_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20109_ _01921_ _01913_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__xor2_2
X_13980_ _06667_ _06678_ _06681_ VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_244_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21089_ net1097 _05328_ _02850_ _02851_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_233_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1054 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12931_ top_inst.grid_inst.data_path_wires\[1\]\[0\] VGND VGND VPWR VPWR _05734_
+ sky130_fd_sc_hd__buf_4
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[12\] _05634_ _05667_
+ _05668_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_69_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _08197_ _08267_ VGND VGND VPWR VPWR _08268_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _07064_ VGND VGND VPWR VPWR _07292_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11813_ net393 _04903_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__or2_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _08159_ _08200_ VGND VGND VPWR VPWR _08201_ sky130_fd_sc_hd__nand2_2
X_12793_ _05599_ _05600_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _09861_ _09862_ VGND VGND VPWR VPWR _09863_ sky130_fd_sc_hd__nand2_1
X_14532_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[6\] _07224_ _06701_
+ VGND VGND VPWR VPWR _07225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11744_ top_inst.axis_out_inst.out_buff_data\[121\] _04865_ VGND VGND VPWR VPWR _04866_
+ sky130_fd_sc_hd__or2_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17251_ _09795_ _09796_ VGND VGND VPWR VPWR _09797_ sky130_fd_sc_hd__xor2_1
XFILLER_0_194_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14463_ _07156_ _07157_ VGND VGND VPWR VPWR _07158_ sky130_fd_sc_hd__nor2_1
XFILLER_0_193_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16202_ _08762_ _08786_ VGND VGND VPWR VPWR _08787_ sky130_fd_sc_hd__nand2_1
X_13414_ top_inst.grid_inst.data_path_wires\[2\]\[1\] VGND VGND VPWR VPWR _06184_
+ sky130_fd_sc_hd__clkbuf_4
X_17182_ _09623_ _09729_ _09730_ VGND VGND VPWR VPWR _09731_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_24_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14394_ _07062_ _07061_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _07093_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16133_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[2\] _07866_ VGND
+ VGND VPWR VPWR _08721_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13345_ _06085_ _06118_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16064_ _08667_ _08140_ VGND VGND VPWR VPWR _08668_ sky130_fd_sc_hd__or2_1
X_13276_ _05980_ _06016_ _06051_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__nor3_1
XFILLER_0_161_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15015_ _07659_ _07660_ VGND VGND VPWR VPWR _07668_ sky130_fd_sc_hd__or2b_1
XFILLER_0_161_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12227_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[5\] _05143_
+ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19823_ _01621_ _01645_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__and2_1
XFILLER_0_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12158_ net310 _05102_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__or2_1
XFILLER_0_208_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19754_ _01569_ _01580_ _01581_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__nand3_1
X_16966_ net204 net201 _09520_ VGND VGND VPWR VPWR _09521_ sky130_fd_sc_hd__nand3_4
X_12089_ net1100 _05063_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18705_ _11145_ _11133_ VGND VGND VPWR VPWR _11146_ sky130_fd_sc_hd__or2_1
X_15917_ _08516_ _08492_ _08527_ VGND VGND VPWR VPWR _08528_ sky130_fd_sc_hd__a21o_1
XFILLER_0_223_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19685_ _01384_ _01429_ _01467_ _01511_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__or4b_4
X_16897_ _09409_ _09449_ _09452_ VGND VGND VPWR VPWR _09453_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_182_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18636_ _11074_ _11093_ _11094_ _05309_ _04861_ VGND VGND VPWR VPWR _11095_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_95_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _08458_ _08460_ VGND VGND VPWR VPWR _08461_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18567_ _10986_ _10988_ VGND VGND VPWR VPWR _11028_ sky130_fd_sc_hd__or2b_1
XFILLER_0_86_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15779_ _08349_ _08393_ VGND VGND VPWR VPWR _08394_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17518_ _10042_ _09199_ VGND VGND VPWR VPWR _10043_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18498_ _10881_ _10916_ _10955_ _10959_ _10954_ VGND VGND VPWR VPWR _10960_ sky130_fd_sc_hd__a32o_1
XFILLER_0_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17449_ _09947_ VGND VGND VPWR VPWR _09986_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_928 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20460_ _02242_ _02243_ _02241_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_244_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19119_ _11536_ _11537_ VGND VGND VPWR VPWR _11538_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20391_ _02144_ _02145_ _02146_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22130_ _03779_ _03784_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__or2b_1
XFILLER_0_70_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22061_ top_inst.deskew_buff_inst.col_input\[99\] _05730_ VGND VGND VPWR VPWR _03755_
+ sky130_fd_sc_hd__and2_1
XTAP_6609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21012_ _02777_ _02778_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22963_ top_inst.skew_buff_inst.row\[1\].output_reg\[1\] _04570_ VGND VGND VPWR VPWR
+ _04571_ sky130_fd_sc_hd__or2_1
XFILLER_0_242_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_94_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_16
X_21914_ _03576_ _03630_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__or2_1
XFILLER_0_218_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22894_ net296 _04522_ _04531_ _04524_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24633_ clknet_leaf_24_clk net628 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[109\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21845_ _03539_ _03565_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24564_ clknet_leaf_134_clk _01097_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dfxtp_4
X_21776_ _03490_ _03498_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23515_ clknet_leaf_137_clk _00048_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20727_ _02502_ _02504_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24495_ clknet_leaf_125_clk _01028_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_184_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23446_ net834 _04840_ _04845_ _04844_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20658_ _02020_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[0\] _02003_
+ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23377_ net460 _04804_ _04807_ _04808_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20589_ _02366_ _02370_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__xnor2_1
X_13130_ _05865_ _05909_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__xnor2_1
X_22328_ _03980_ _03979_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__or2b_1
XFILLER_0_108_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13061_ _05840_ _05842_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__xnor2_1
X_22259_ top_inst.grid_inst.data_path_wires\[18\]\[6\] top_inst.grid_inst.data_path_wires\[18\]\[5\]
+ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1097 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12012_ _04994_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__buf_2
XFILLER_0_218_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16820_ _09360_ _09377_ _09186_ _09191_ VGND VGND VPWR VPWR _09378_ sky130_fd_sc_hd__or4b_4
XFILLER_0_205_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16751_ _09302_ _09303_ _09310_ VGND VGND VPWR VPWR _09311_ sky130_fd_sc_hd__and3_1
XFILLER_0_219_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13963_ _06680_ _06681_ _06682_ VGND VGND VPWR VPWR _06683_ sky130_fd_sc_hd__a21o_1
XFILLER_0_221_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_85_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_216_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15702_ top_inst.grid_inst.data_path_wires\[7\]\[4\] top_inst.grid_inst.data_path_wires\[7\]\[3\]
+ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _08318_ sky130_fd_sc_hd__nand4_2
X_12914_ _05691_ _05695_ _05717_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__a21o_1
X_19470_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[7\] _01303_ VGND
+ VGND VPWR VPWR _01304_ sky130_fd_sc_hd__xor2_2
X_16682_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[2\] _08066_ _09243_
+ _09244_ VGND VGND VPWR VPWR _09245_ sky130_fd_sc_hd__a22o_1
X_13894_ _06628_ _06620_ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18421_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[9\] _10793_ _10840_
+ VGND VGND VPWR VPWR _10885_ sky130_fd_sc_hd__a21o_1
XFILLER_0_243_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12845_ _05638_ _05610_ _05650_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__nand3_1
XFILLER_0_198_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15633_ top_inst.grid_inst.data_path_wires\[7\]\[5\] top_inst.grid_inst.data_path_wires\[7\]\[4\]
+ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[1\] _08154_ VGND VGND
+ VPWR VPWR _08251_ sky130_fd_sc_hd__nand4_1
XFILLER_0_150_1013 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _10788_ _10817_ VGND VGND VPWR VPWR _10818_ sky130_fd_sc_hd__xnor2_1
X_12776_ _05579_ _05580_ _05584_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__nand3_1
XFILLER_0_115_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15564_ _08139_ _08137_ _08157_ _08155_ VGND VGND VPWR VPWR _08185_ sky130_fd_sc_hd__nand4_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17303_ _09819_ _09846_ VGND VGND VPWR VPWR _09847_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14515_ _07202_ _07203_ _07206_ VGND VGND VPWR VPWR _07208_ sky130_fd_sc_hd__a21o_1
X_15495_ _06848_ _08133_ _08134_ _07643_ VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__o211a_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18283_ _10716_ _10722_ VGND VGND VPWR VPWR _10750_ sky130_fd_sc_hd__or2b_1
XFILLER_0_189_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17234_ _09777_ _09780_ VGND VGND VPWR VPWR _09781_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14446_ _07138_ _07139_ _07127_ VGND VGND VPWR VPWR _07141_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14377_ _07079_ _07075_ VGND VGND VPWR VPWR _07080_ sky130_fd_sc_hd__or2_1
X_17165_ _09698_ _09714_ VGND VGND VPWR VPWR _09715_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold907 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[12\] VGND VGND
+ VPWR VPWR net1089 sky130_fd_sc_hd__dlygate4sd3_1
X_13328_ _06101_ _06102_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__xnor2_1
X_16116_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[1\] _08703_ _08704_
+ VGND VGND VPWR VPWR _08705_ sky130_fd_sc_hd__nand3_1
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold918 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[10\] VGND
+ VGND VPWR VPWR net1100 sky130_fd_sc_hd__dlygate4sd3_1
X_17096_ _09645_ _09646_ _09634_ VGND VGND VPWR VPWR _09648_ sky130_fd_sc_hd__a21o_1
Xhold929 top_inst.axis_in_inst.inbuf_bus\[19\] VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_724 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13259_ _06032_ _06034_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__and2_1
X_16047_ _08532_ _08630_ _08653_ VGND VGND VPWR VPWR _08654_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_228_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19806_ _01611_ _01610_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17998_ _10056_ _10499_ _10460_ _10500_ VGND VGND VPWR VPWR _10501_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_97_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19737_ _01526_ _01530_ _01564_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__a21o_1
X_16949_ _09502_ _09503_ VGND VGND VPWR VPWR _09504_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_237_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_76_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_189_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19668_ _01495_ _01496_ _01488_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18619_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[15\] _10923_ VGND
+ VGND VPWR VPWR _11078_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_189_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19599_ net464 _01386_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__or2_1
XFILLER_0_176_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21630_ _03349_ _03350_ _03358_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__or3_1
XFILLER_0_192_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21561_ _03253_ _03291_ _03292_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__a21o_1
XFILLER_0_191_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23300_ net142 _04753_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20512_ _02240_ _02247_ _02246_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_51_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24280_ clknet_leaf_11_clk _00813_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[17\]\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21492_ _03223_ _03225_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__xor2_2
XFILLER_0_172_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23231_ net109 _04714_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20443_ _01990_ _02227_ _02189_ _02190_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_144_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23162_ _04684_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__clkbuf_4
X_20374_ _02157_ _02158_ _02159_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_141_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22113_ _03311_ _03804_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23093_ net580 _10541_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__nand2_1
XTAP_6406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22044_ _03729_ _03730_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__nand2_1
XTAP_6439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23995_ clknet_leaf_79_clk _00528_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_243_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_242_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22946_ top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[2\] _04557_ VGND
+ VGND VPWR VPWR _04561_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22877_ net809 _04509_ _04521_ _04511_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12630_ _05432_ _05433_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__and2b_1
XFILLER_0_210_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24616_ clknet_leaf_31_clk _01149_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_156_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21828_ _03469_ _03546_ _03548_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__a21o_1
XFILLER_0_183_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_1388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12561_ _05375_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24547_ clknet_leaf_100_clk _01080_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_66_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21759_ _03460_ _03483_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14300_ _07007_ _07009_ VGND VGND VPWR VPWR _07010_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15280_ _07624_ _07631_ _07877_ _07878_ VGND VGND VPWR VPWR _07926_ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24478_ clknet_leaf_37_clk _01011_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12492_ _05310_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__buf_8
XFILLER_0_0_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14231_ _06941_ _06942_ VGND VGND VPWR VPWR _06943_ sky130_fd_sc_hd__nor2_1
XFILLER_0_227_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23429_ top_inst.axis_out_inst.out_buff_data\[103\] _04835_ VGND VGND VPWR VPWR _04836_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_62_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire167 _11129_ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_4
XFILLER_0_180_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14162_ _06777_ _06779_ _06826_ VGND VGND VPWR VPWR _06876_ sky130_fd_sc_hd__and3_1
XFILLER_0_151_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13113_ _05891_ _05892_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14093_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[3\]\[2\]
+ _06806_ VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__and3_1
X_18970_ _11390_ _11391_ VGND VGND VPWR VPWR _11392_ sky130_fd_sc_hd__nor2_1
XFILLER_0_237_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13044_ _05824_ _05825_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__nand2_1
X_17921_ _10379_ _10381_ VGND VGND VPWR VPWR _10426_ sky130_fd_sc_hd__nor2_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17852_ _10357_ _10358_ VGND VGND VPWR VPWR _10359_ sky130_fd_sc_hd__and2_1
XFILLER_0_234_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16803_ _09360_ VGND VGND VPWR VPWR _09361_ sky130_fd_sc_hd__buf_2
XFILLER_0_79_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17783_ _10244_ _10253_ VGND VGND VPWR VPWR _10291_ sky130_fd_sc_hd__or2b_1
Xclkbuf_leaf_58_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_16
X_14995_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[1\] _07648_ _07649_
+ VGND VGND VPWR VPWR _07650_ sky130_fd_sc_hd__nand3_2
X_19522_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[8\] _01354_ VGND
+ VGND VPWR VPWR _01355_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_221_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16734_ _09262_ _09289_ VGND VGND VPWR VPWR _09294_ sky130_fd_sc_hd__nor2_1
X_13946_ _06662_ _06663_ _06664_ _06665_ VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__nand4_2
XFILLER_0_72_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19453_ net237 _01286_ _01247_ _01260_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16665_ _09226_ _09227_ _09222_ VGND VGND VPWR VPWR _09229_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_158_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_1287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13877_ _06609_ _06610_ _06615_ _05313_ VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_57_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18404_ _10796_ _10813_ _10868_ VGND VGND VPWR VPWR _10869_ sky130_fd_sc_hd__a21oi_1
X_15616_ _08233_ _08234_ VGND VGND VPWR VPWR _08235_ sky130_fd_sc_hd__nor2_1
X_12828_ _05626_ _05627_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__or2b_1
X_19384_ _01218_ _01219_ _01220_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__or3b_4
XFILLER_0_189_1020 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16596_ _09165_ _09167_ _09168_ _09170_ _05313_ VGND VGND VPWR VPWR _09171_ sky130_fd_sc_hd__o311a_1
XFILLER_0_201_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18335_ _10799_ _10800_ VGND VGND VPWR VPWR _10801_ sky130_fd_sc_hd__nand2_1
XFILLER_0_210_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15547_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[7\] _07641_ VGND
+ VGND VPWR VPWR _08171_ sky130_fd_sc_hd__or2_1
X_12759_ _05447_ _05449_ _05287_ _05567_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__or4_1
XFILLER_0_173_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18266_ _10724_ _10733_ VGND VGND VPWR VPWR _10734_ sky130_fd_sc_hd__xor2_1
XFILLER_0_155_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15478_ _08094_ _08095_ _08092_ VGND VGND VPWR VPWR _08119_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17217_ _09741_ _09744_ _09764_ VGND VGND VPWR VPWR _09765_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_141_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14429_ _07123_ _07124_ VGND VGND VPWR VPWR _07125_ sky130_fd_sc_hd__or2b_1
XFILLER_0_181_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18197_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[4\] _10666_ VGND
+ VGND VPWR VPWR _10667_ sky130_fd_sc_hd__xor2_2
XFILLER_0_141_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17148_ _09688_ _09666_ VGND VGND VPWR VPWR _09698_ sky130_fd_sc_hd__and2b_1
XFILLER_0_130_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold704 top_inst.deskew_buff_inst.col_input\[84\] VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold715 top_inst.deskew_buff_inst.col_input\[74\] VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold726 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[21\] VGND
+ VGND VPWR VPWR net908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold737 top_inst.deskew_buff_inst.col_input\[57\] VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold748 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[0\] VGND
+ VGND VPWR VPWR net930 sky130_fd_sc_hd__dlygate4sd3_1
X_17079_ _09419_ VGND VGND VPWR VPWR _09631_ sky130_fd_sc_hd__clkbuf_8
Xhold759 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[12\] VGND
+ VGND VPWR VPWR net941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20090_ _01901_ _01902_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22800_ _04432_ _04431_ _04448_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23780_ clknet_leaf_65_clk _00313_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20992_ net919 _02491_ _02758_ _02759_ _01863_ VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__o221a_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22731_ _04401_ _04402_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__nor2_1
XFILLER_0_211_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22662_ _04319_ _04336_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24401_ clknet_leaf_57_clk net397 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].output_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21613_ _03339_ _03342_ _10831_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__o21a_1
XFILLER_0_164_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22593_ _04261_ _04270_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24332_ clknet_leaf_5_clk _00865_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_62_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21544_ _03239_ _03271_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24263_ clknet_leaf_110_clk _00796_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21475_ _03168_ _03208_ VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__nor2_2
XFILLER_0_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23214_ net101 _04714_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20426_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[7\] _02210_ _02211_
+ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24194_ clknet_leaf_117_clk _00727_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23145_ net69 _04672_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__or2_1
X_20357_ _01989_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[5\] VGND
+ VGND VPWR VPWR _02144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_219_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23076_ top_inst.axis_in_inst.inbuf_bus\[25\] _04629_ VGND VGND VPWR VPWR _04636_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_235_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20288_ _01989_ _01986_ _02013_ _02011_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__and4_1
XTAP_5502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22027_ _03715_ _03720_ _03721_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__nand3_1
XTAP_6269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold75 _00162_ VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold86 top_inst.deskew_buff_inst.col_input\[50\] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ _06537_ _06542_ VGND VGND VPWR VPWR _06543_ sky130_fd_sc_hd__xnor2_1
Xhold97 _00118_ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_243_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14780_ _07456_ _07457_ _07466_ VGND VGND VPWR VPWR _07467_ sky130_fd_sc_hd__a21o_1
XFILLER_0_199_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11992_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[0\] _05010_
+ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__or2_1
XTAP_4889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23978_ clknet_leaf_87_clk _00511_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_216_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13731_ _06436_ _06438_ _06475_ VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__o21a_1
X_22929_ net662 _04543_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__or2_1
XFILLER_0_230_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16450_ _08978_ _08977_ VGND VGND VPWR VPWR _09029_ sky130_fd_sc_hd__or2b_1
XFILLER_0_116_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13662_ _06399_ _06401_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15401_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[13\] _07924_ VGND
+ VGND VPWR VPWR _08044_ sky130_fd_sc_hd__xnor2_1
X_12613_ _05424_ _05425_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_1196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16381_ _08697_ _08671_ _08669_ _08876_ VGND VGND VPWR VPWR _08961_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_137_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13593_ _06299_ _06301_ VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__nand2_1
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18120_ _10600_ _10057_ VGND VGND VPWR VPWR _10601_ sky130_fd_sc_hd__or2_1
X_12544_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[1\] _05286_ _05291_
+ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _05359_ sky130_fd_sc_hd__a22oi_1
X_15332_ _07923_ _07929_ _07921_ VGND VGND VPWR VPWR _07977_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18051_ _10547_ _10551_ VGND VGND VPWR VPWR _10552_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12475_ _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__buf_4
X_15263_ _07613_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[7\] _07640_
+ _07615_ VGND VGND VPWR VPWR _07909_ sky130_fd_sc_hd__and4b_1
XFILLER_0_48_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17002_ _09361_ _09205_ _09209_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _09556_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_152_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14214_ _06652_ top_inst.grid_inst.data_path_wires\[3\]\[5\] _06925_ VGND VGND VPWR
+ VPWR _06926_ sky130_fd_sc_hd__a21oi_1
X_15194_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[1\] _07626_ top_inst.grid_inst.data_path_wires\[6\]\[7\]
+ VGND VGND VPWR VPWR _07842_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_6 _08265_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_227_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14145_ _06857_ _06858_ VGND VGND VPWR VPWR _06859_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_240_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_238_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14076_ _06782_ _06791_ VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__xor2_2
XFILLER_0_123_1254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18953_ _11288_ _11327_ VGND VGND VPWR VPWR _11376_ sky130_fd_sc_hd__nor2_1
XFILLER_0_238_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13027_ _05741_ _05761_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__nand2_1
X_17904_ _10387_ _10389_ VGND VGND VPWR VPWR _10409_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18884_ _11274_ _11279_ VGND VGND VPWR VPWR _11308_ sky130_fd_sc_hd__and2_1
XTAP_6770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17835_ _10340_ _10341_ VGND VGND VPWR VPWR _10342_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer18 _09464_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17766_ _10271_ _10273_ _08265_ VGND VGND VPWR VPWR _10275_ sky130_fd_sc_hd__o21a_1
Xrebuffer29 _05266_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__buf_4
XFILLER_0_178_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14978_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _07637_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19505_ _01335_ _01337_ _01287_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16717_ _09255_ _09276_ _09277_ VGND VGND VPWR VPWR _09278_ sky130_fd_sc_hd__or3_4
XFILLER_0_77_806 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13929_ _06632_ _06647_ _06653_ _06639_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__o211a_1
X_17697_ _10035_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[2\] _10205_
+ _10206_ VGND VGND VPWR VPWR _10207_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1035 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19436_ _11697_ _11693_ _11687_ _11692_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__nand4_2
X_16648_ _09214_ VGND VGND VPWR VPWR _09215_ sky130_fd_sc_hd__buf_2
XFILLER_0_159_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19367_ _11683_ _11678_ net234 _11696_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__nand4_1
XFILLER_0_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16579_ _09055_ _09153_ VGND VGND VPWR VPWR _09154_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18318_ _10783_ _10784_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[7\]
+ _07816_ VGND VGND VPWR VPWR _10785_ sky130_fd_sc_hd__a2bb2o_1
X_19298_ _11697_ _11689_ VGND VGND VPWR VPWR _11698_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18249_ _10604_ _10686_ _10688_ _10685_ VGND VGND VPWR VPWR _10717_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_199_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21260_ _02889_ _02967_ _02969_ _02966_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_128_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold501 _00066_ VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold512 top_inst.axis_out_inst.out_buff_data\[90\] VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 top_inst.axis_out_inst.out_buff_data\[76\] VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__dlygate4sd3_1
X_20211_ _01990_ _11163_ _02010_ _02006_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold534 _00918_ VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold545 top_inst.axis_out_inst.out_buff_data\[75\] VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__dlygate4sd3_1
X_21191_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[2\] _02911_ _02912_
+ VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_141_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold556 _00103_ VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold567 top_inst.axis_out_inst.out_buff_data\[28\] VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20142_ _01563_ _01952_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold578 top_inst.deskew_buff_inst.col_input\[33\] VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[6\] VGND VGND
+ VPWR VPWR net771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_244_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20073_ _05887_ _01885_ _01886_ _01887_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__a31o_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23901_ clknet_4_13__leaf_clk _00434_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23832_ clknet_leaf_93_clk _00365_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23763_ clknet_leaf_66_clk _00296_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_20975_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[25\] _02470_ VGND
+ VGND VPWR VPWR _02743_ sky130_fd_sc_hd__or2_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22714_ _04369_ _04372_ _04371_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23694_ clknet_leaf_119_clk _00227_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22645_ _04319_ _04320_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22576_ _04205_ _04208_ _04233_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24315_ clknet_leaf_1_clk _00848_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[90\]
+ sky130_fd_sc_hd__dfxtp_1
X_21527_ _03257_ _03259_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__xor2_2
XFILLER_0_106_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24246_ clknet_leaf_108_clk _00779_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_12260_ net678 _05156_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__or2_1
X_21458_ _03190_ _03192_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__nand2_1
XFILLER_0_224_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_1216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20409_ top_inst.grid_inst.data_path_wires\[16\]\[6\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[1\]
+ _02192_ _02193_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__a22o_1
X_24177_ clknet_leaf_29_clk _00710_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_12191_ _05044_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__clkbuf_4
X_21389_ _03084_ _03087_ _03085_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_102_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23128_ net121 _04659_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__or2_1
Xoutput43 net43 VGND VGND VPWR VPWR output_tdata[104] sky130_fd_sc_hd__clkbuf_4
Xoutput54 net54 VGND VGND VPWR VPWR output_tdata[114] sky130_fd_sc_hd__clkbuf_4
XTAP_6011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput65 net65 VGND VGND VPWR VPWR output_tdata[124] sky130_fd_sc_hd__clkbuf_4
XTAP_6022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput76 net76 VGND VGND VPWR VPWR output_tdata[19] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_235_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput87 net87 VGND VGND VPWR VPWR output_tdata[29] sky130_fd_sc_hd__clkbuf_4
XTAP_6055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23059_ net994 _04616_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__or2_1
XTAP_5310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15950_ _08150_ _08353_ _08558_ VGND VGND VPWR VPWR _08560_ sky130_fd_sc_hd__nor3_1
Xoutput98 net98 VGND VGND VPWR VPWR output_tdata[39] sky130_fd_sc_hd__buf_2
XTAP_5321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14901_ _07563_ _07583_ VGND VGND VPWR VPWR _07584_ sky130_fd_sc_hd__xnor2_1
XTAP_6088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15881_ _08484_ _08491_ VGND VGND VPWR VPWR _08493_ sky130_fd_sc_hd__or2_1
XFILLER_0_208_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ _10128_ _10131_ VGND VGND VPWR VPWR _10132_ sky130_fd_sc_hd__xor2_2
X_14832_ _07483_ _07480_ _07517_ VGND VGND VPWR VPWR _07518_ sky130_fd_sc_hd__a21oi_1
XTAP_5398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1068 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_975 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _10064_ _10065_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[1\]
+ VGND VGND VPWR VPWR _10067_ sky130_fd_sc_hd__a21o_1
X_14763_ _07328_ _07413_ _07412_ VGND VGND VPWR VPWR _07450_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_187_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ net791 _04990_ _05000_ _04995_ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ net1008 _05403_ VGND VGND VPWR VPWR _09079_ sky130_fd_sc_hd__nand2_1
XTAP_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13714_ _06195_ _06210_ _06208_ top_inst.grid_inst.data_path_wires\[2\]\[7\] VGND
+ VGND VPWR VPWR _06459_ sky130_fd_sc_hd__a22oi_1
X_17482_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[25\] _10015_ _09418_
+ VGND VGND VPWR VPWR _10016_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14694_ _07381_ _07382_ VGND VGND VPWR VPWR _07383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19221_ _11635_ _11636_ VGND VGND VPWR VPWR _11637_ sky130_fd_sc_hd__and2_1
X_16433_ _09010_ _09011_ VGND VGND VPWR VPWR _09012_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_195_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13645_ _06389_ _06391_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19152_ _11557_ _11529_ _11568_ VGND VGND VPWR VPWR _11570_ sky130_fd_sc_hd__nand3_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16364_ _08891_ _08889_ VGND VGND VPWR VPWR _08945_ sky130_fd_sc_hd__and2b_1
XFILLER_0_13_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13576_ _06322_ _06324_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[6\]
+ _05327_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_171_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18103_ _10032_ _10584_ _10588_ _10448_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15315_ _07958_ _07959_ VGND VGND VPWR VPWR _07960_ sky130_fd_sc_hd__and2b_1
X_12527_ _05280_ _05283_ _05342_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__nand3_1
X_19083_ _11460_ _11463_ _11501_ _10957_ VGND VGND VPWR VPWR _11503_ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16295_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[8\]\[2\]
+ top_inst.grid_inst.data_path_wires\[8\]\[1\] _08876_ VGND VGND VPWR VPWR _08877_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18034_ _10534_ _10535_ VGND VGND VPWR VPWR _10536_ sky130_fd_sc_hd__or2_1
X_15246_ _07886_ _07892_ VGND VGND VPWR VPWR _07893_ sky130_fd_sc_hd__xnor2_1
X_12458_ _05282_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__buf_2
XFILLER_0_140_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15177_ top_inst.grid_inst.data_path_wires\[6\]\[2\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[6\]
+ _07824_ top_inst.grid_inst.data_path_wires\[6\]\[1\] VGND VGND VPWR VPWR _07825_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12389_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[11\] _05235_
+ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14128_ _06800_ _06798_ VGND VGND VPWR VPWR _06843_ sky130_fd_sc_hd__or2b_1
X_19985_ _01561_ _01802_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14059_ _06741_ _06774_ VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__xor2_2
X_18936_ _11273_ _11318_ VGND VGND VPWR VPWR _11359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_1152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1027 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18867_ _11290_ _11291_ VGND VGND VPWR VPWR _11292_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17818_ _10310_ _10312_ VGND VGND VPWR VPWR _10325_ sky130_fd_sc_hd__or2_1
X_18798_ _11203_ _11205_ VGND VGND VPWR VPWR _11225_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17749_ _10239_ _10257_ VGND VGND VPWR VPWR _10258_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20760_ _02455_ _02536_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19419_ _01250_ _01251_ _01253_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20691_ _02467_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__buf_2
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22430_ _04112_ _04113_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__xor2_1
XFILLER_0_174_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22361_ _04012_ _04008_ _04046_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24100_ clknet_leaf_15_clk _00633_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_116_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21312_ top_inst.grid_inst.data_path_wires\[17\]\[2\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[5\]
+ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22292_ _03695_ _03703_ _03946_ _03947_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24031_ clknet_leaf_48_clk _00564_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold320 _00152_ VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__dlygate4sd3_1
X_21243_ _02948_ _02949_ _02982_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold331 top_inst.axis_out_inst.out_buff_data\[44\] VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold342 top_inst.deskew_buff_inst.col_input\[88\] VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[11\] VGND
+ VGND VPWR VPWR net535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[7\] VGND
+ VGND VPWR VPWR net546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 top_inst.axis_out_inst.out_buff_data\[95\] VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__dlygate4sd3_1
X_21174_ _02910_ _02916_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__or2_1
XFILLER_0_159_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold386 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[8\] VGND
+ VGND VPWR VPWR net568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 _00903_ VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_244_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_217_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20125_ _01563_ _01935_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_244_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20056_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[25\] _01761_ _01762_
+ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__a21o_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23815_ clknet_leaf_72_clk _00348_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11760_ net564 _04860_ _04878_ _04875_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__o211a_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20958_ _02725_ _02726_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__and2_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23746_ clknet_leaf_122_clk _00279_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20889_ net782 _02638_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__or2_1
X_23677_ clknet_leaf_116_clk net421 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13430_ top_inst.grid_inst.data_path_wires\[2\]\[6\] VGND VGND VPWR VPWR _06195_
+ sky130_fd_sc_hd__buf_2
X_22628_ net533 _09804_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13361_ _06065_ _06103_ _06134_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22559_ _04199_ _04237_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15100_ _07615_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[2\] _07748_
+ _07749_ VGND VGND VPWR VPWR _07750_ sky130_fd_sc_hd__a22o_1
Xrebuffer9 net190 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__buf_1
X_12312_ net807 _05183_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16080_ top_inst.grid_inst.data_path_wires\[8\]\[7\] VGND VGND VPWR VPWR _08679_
+ sky130_fd_sc_hd__clkbuf_4
X_13292_ _06063_ _06067_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15031_ _07667_ _07682_ _07683_ VGND VGND VPWR VPWR _07684_ sky130_fd_sc_hd__or3_1
X_12243_ net826 _05151_ _05153_ _05141_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__o211a_1
X_24229_ clknet_leaf_113_clk _00762_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[16\]\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_224_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12174_ _04994_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19770_ _01565_ _01587_ _01585_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16982_ _05399_ _09536_ VGND VGND VPWR VPWR _09537_ sky130_fd_sc_hd__nor2_1
X_18721_ _11156_ _11150_ VGND VGND VPWR VPWR _11157_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15933_ _08505_ _08507_ VGND VGND VPWR VPWR _08544_ sky130_fd_sc_hd__or2b_1
XFILLER_0_120_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18652_ _11087_ _11076_ VGND VGND VPWR VPWR _11110_ sky130_fd_sc_hd__and2b_1
XTAP_5195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[11\] VGND VGND
+ VPWR VPWR _08476_ sky130_fd_sc_hd__inv_2
XTAP_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ _10052_ _10088_ _10115_ VGND VGND VPWR VPWR _10116_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_235_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14815_ _07495_ _07500_ VGND VGND VPWR VPWR _07501_ sky130_fd_sc_hd__xnor2_1
XTAP_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18583_ _11011_ _11026_ _11024_ VGND VGND VPWR VPWR _11043_ sky130_fd_sc_hd__o21a_1
XTAP_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15795_ top_inst.grid_inst.data_path_wires\[7\]\[7\] _08159_ VGND VGND VPWR VPWR
+ _08409_ sky130_fd_sc_hd__nand2_4
XFILLER_0_192_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_235_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17534_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _10054_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_114_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14746_ _07404_ _07433_ VGND VGND VPWR VPWR _07434_ sky130_fd_sc_hd__xor2_1
XTAP_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11958_ _04911_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17465_ _09919_ _09957_ _09976_ VGND VGND VPWR VPWR _10001_ sky130_fd_sc_hd__or3_1
XFILLER_0_129_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14677_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[10\] _07281_ VGND
+ VGND VPWR VPWR _07366_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11889_ _04911_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__clkbuf_4
X_19204_ _11610_ _11613_ VGND VGND VPWR VPWR _11620_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16416_ _08992_ _08994_ _08265_ VGND VGND VPWR VPWR _08996_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13628_ top_inst.grid_inst.data_path_wires\[2\]\[4\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[2\]\[5\]
+ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17396_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[25\] _09628_ _09629_
+ VGND VGND VPWR VPWR _09935_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_131_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19135_ _11514_ _11552_ VGND VGND VPWR VPWR _11553_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16347_ _08673_ _08693_ _08690_ _08676_ VGND VGND VPWR VPWR _08928_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13559_ _06306_ _06307_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19066_ _11442_ _11444_ _11443_ VGND VGND VPWR VPWR _11486_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_89_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16278_ _08819_ _08820_ VGND VGND VPWR VPWR _08861_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_242_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18017_ _10479_ _10515_ VGND VGND VPWR VPWR _10519_ sky130_fd_sc_hd__or2b_1
XFILLER_0_125_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15229_ _07874_ _07875_ VGND VGND VPWR VPWR _07876_ sky130_fd_sc_hd__xor2_1
XFILLER_0_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19968_ _01760_ _01771_ _01784_ _01743_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__a22oi_2
X_18919_ _11337_ _11341_ VGND VGND VPWR VPWR _11342_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19899_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[18\] _01395_ _01396_
+ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__a21o_2
XFILLER_0_207_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21930_ _03646_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__inv_2
XFILLER_0_222_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21861_ _03580_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23600_ clknet_leaf_103_clk net560 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20812_ _02556_ _02572_ _02585_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__and3_1
XFILLER_0_195_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24580_ clknet_leaf_142_clk _01113_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dfxtp_4
X_21792_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[21\] _03421_ _03422_
+ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_38_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_212_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23531_ clknet_leaf_142_clk _00064_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20743_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[16\] _02470_ VGND
+ VGND VPWR VPWR _02520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23462_ net884 _04859_ _04853_ _04844_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20674_ _01819_ _02452_ _02453_ _02035_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22413_ _04094_ _04096_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__and2_1
XFILLER_0_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23393_ net739 _04804_ _04816_ _04808_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22344_ _04026_ _04029_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22275_ _03960_ _03962_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24014_ clknet_leaf_48_clk _00547_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_83_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold150 _01022_ VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__dlygate4sd3_1
X_21226_ _02868_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[2\] VGND
+ VGND VPWR VPWR _02966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold161 top_inst.deskew_buff_inst.col_input\[3\] VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 top_inst.valid_pipe\[5\] VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold183 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[23\] VGND
+ VGND VPWR VPWR net365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _00196_ VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21157_ net454 _01735_ _02901_ _02880_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__o211a_1
XFILLER_0_244_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20108_ _01916_ _01920_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__xor2_2
XFILLER_0_176_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21088_ _02840_ _02847_ _05406_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_226_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12930_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[15\] _05314_ _05733_
+ _05308_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_1066 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20039_ _01853_ _01854_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__nand2_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12861_ _05635_ _05629_ _05666_ _05633_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__a31o_1
XFILLER_0_198_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14600_ _07241_ _07242_ _07065_ _07290_ VGND VGND VPWR VPWR _07291_ sky130_fd_sc_hd__or4_4
XFILLER_0_154_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11812_ net800 _04898_ _04907_ _04902_ VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__o211a_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15580_ top_inst.grid_inst.data_path_wires\[7\]\[1\] top_inst.grid_inst.data_path_wires\[7\]\[0\]
+ _08161_ VGND VGND VPWR VPWR _08200_ sky130_fd_sc_hd__and3_1
X_12792_ _05298_ _05301_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14531_ _07221_ _07223_ VGND VGND VPWR VPWR _07224_ sky130_fd_sc_hd__xor2_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _04864_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__buf_4
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23729_ clknet_leaf_121_clk _00262_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17250_ _09726_ _09774_ VGND VGND VPWR VPWR _09796_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14462_ net173 _07112_ _07131_ _07130_ VGND VGND VPWR VPWR _07157_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16201_ _08783_ _08785_ VGND VGND VPWR VPWR _08786_ sky130_fd_sc_hd__xnor2_1
X_13413_ _05734_ _05256_ _06182_ _06183_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__o211a_1
X_17181_ _09588_ _09459_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[16\]
+ VGND VGND VPWR VPWR _09730_ sky130_fd_sc_hd__a21o_1
XFILLER_0_180_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14393_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[7\] _05276_ _07091_
+ _07092_ VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16132_ _08708_ _08719_ VGND VGND VPWR VPWR _08720_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_181_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13344_ _06116_ _06117_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16063_ top_inst.grid_inst.data_path_wires\[8\]\[2\] VGND VGND VPWR VPWR _08667_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13275_ _05765_ _05763_ _05753_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15014_ _07653_ _07664_ VGND VGND VPWR VPWR _07667_ sky130_fd_sc_hd__or2b_1
X_12226_ net355 _05137_ _05144_ _05141_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__o211a_1
XFILLER_0_241_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19822_ net1093 _01202_ _01646_ _01647_ _11228_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__o221a_1
X_12157_ net418 _05097_ _05104_ _05101_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16965_ _09469_ _09477_ _09476_ VGND VGND VPWR VPWR _09520_ sky130_fd_sc_hd__a21bo_2
X_19753_ _01577_ _01578_ _01579_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__a21o_1
X_12088_ net577 _05058_ _05065_ _05062_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18704_ top_inst.grid_inst.data_path_wires\[13\]\[6\] VGND VGND VPWR VPWR _11145_
+ sky130_fd_sc_hd__buf_2
X_15916_ _08525_ _08526_ VGND VGND VPWR VPWR _08527_ sky130_fd_sc_hd__nand2_1
X_19684_ net1092 _01202_ _01512_ _01513_ _11228_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__o221a_1
X_16896_ _09447_ _09448_ VGND VGND VPWR VPWR _09452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18635_ _11074_ _11093_ VGND VGND VPWR VPWR _11094_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ _08414_ _08420_ _08459_ VGND VGND VPWR VPWR _08460_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_177_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18566_ _11011_ _11026_ VGND VGND VPWR VPWR _11027_ sky130_fd_sc_hd__xor2_2
XTAP_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15778_ _08391_ _08392_ VGND VGND VPWR VPWR _08393_ sky130_fd_sc_hd__and2_1
XFILLER_0_176_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17517_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _10042_ sky130_fd_sc_hd__clkbuf_4
X_14729_ _07241_ _07242_ _07078_ _07416_ VGND VGND VPWR VPWR _07417_ sky130_fd_sc_hd__or4_1
XFILLER_0_157_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18497_ _10911_ _10914_ VGND VGND VPWR VPWR _10959_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17448_ _09965_ _09983_ VGND VGND VPWR VPWR _09985_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17379_ _09726_ VGND VGND VPWR VPWR _09919_ sky130_fd_sc_hd__buf_2
XFILLER_0_172_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19118_ _11535_ _11511_ VGND VGND VPWR VPWR _11537_ sky130_fd_sc_hd__or2b_1
XFILLER_0_54_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20390_ _02168_ _02175_ _02171_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19049_ _11340_ VGND VGND VPWR VPWR _11469_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22060_ _03751_ _03752_ _03737_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21011_ _02754_ _02776_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_1088 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22962_ _04863_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__buf_2
XFILLER_0_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21913_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[27\] _03421_ _03422_
+ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_241_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22893_ top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[3\] _04530_ VGND
+ VGND VPWR VPWR _04531_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24632_ clknet_leaf_23_clk net660 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[108\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21844_ _03563_ _03564_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__and2_1
XFILLER_0_214_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24563_ clknet_leaf_137_clk _01096_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dfxtp_4
X_21775_ _03490_ _03498_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23514_ clknet_leaf_137_clk _00047_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_20726_ _02463_ _02476_ _02503_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24494_ clknet_leaf_108_clk _01027_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_147_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23445_ net423 _04835_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20657_ _02365_ _02407_ _02364_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23376_ _04690_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20588_ _02368_ _02369_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22327_ _04003_ _03976_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__or2b_1
XFILLER_0_108_1130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13060_ _05795_ _05816_ _05841_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__o21a_1
X_22258_ top_inst.grid_inst.data_path_wires\[18\]\[5\] top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[18\]\[6\]
+ VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12011_ net577 _05010_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21209_ _02948_ _02949_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__xnor2_2
X_22189_ _03713_ _03878_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_217_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_233_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16750_ _09308_ _09309_ VGND VGND VPWR VPWR _09310_ sky130_fd_sc_hd__nor2_1
X_13962_ _05327_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__buf_6
XFILLER_0_219_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15701_ top_inst.grid_inst.data_path_wires\[7\]\[3\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[7\]\[4\]
+ VGND VGND VPWR VPWR _08317_ sky130_fd_sc_hd__a22o_1
X_12913_ _05691_ _05695_ _05717_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16681_ _09229_ _09242_ _08265_ VGND VGND VPWR VPWR _09244_ sky130_fd_sc_hd__o21a_1
XFILLER_0_216_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13893_ top_inst.grid_inst.data_path_wires\[3\]\[4\] VGND VGND VPWR VPWR _06628_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18420_ _10841_ _10845_ _10843_ VGND VGND VPWR VPWR _10884_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15632_ top_inst.grid_inst.data_path_wires\[7\]\[4\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[1\]
+ _08154_ top_inst.grid_inst.data_path_wires\[7\]\[5\] VGND VGND VPWR VPWR _08250_
+ sky130_fd_sc_hd__a22o_1
X_12844_ _05638_ _05610_ _05650_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _10814_ _10816_ VGND VGND VPWR VPWR _10817_ sky130_fd_sc_hd__xor2_1
X_15563_ _08137_ _08157_ _08155_ _08139_ VGND VGND VPWR VPWR _08184_ sky130_fd_sc_hd__a22o_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12775_ _05582_ _05583_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__and2_1
XFILLER_0_201_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _09844_ _09845_ VGND VGND VPWR VPWR _09846_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14514_ _07202_ _07203_ _07206_ VGND VGND VPWR VPWR _07207_ sky130_fd_sc_hd__nand3_1
XFILLER_0_185_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ _10749_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__clkbuf_1
X_15494_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[16\] _07866_ VGND
+ VGND VPWR VPWR _08134_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17233_ _09778_ _09775_ _09779_ VGND VGND VPWR VPWR _09780_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14445_ _07127_ _07138_ _07139_ VGND VGND VPWR VPWR _07140_ sky130_fd_sc_hd__or3_1
XFILLER_0_181_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17164_ _09712_ _09713_ VGND VGND VPWR VPWR _09714_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14376_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _07079_ sky130_fd_sc_hd__buf_2
XFILLER_0_163_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16115_ _08686_ _08664_ _08683_ _08661_ VGND VGND VPWR VPWR _08704_ sky130_fd_sc_hd__nand4_1
Xhold908 top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[12\] VGND VGND
+ VPWR VPWR net1090 sky130_fd_sc_hd__dlygate4sd3_1
X_13327_ _06063_ _06067_ _06061_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17095_ _09634_ _09645_ _09646_ VGND VGND VPWR VPWR _09647_ sky130_fd_sc_hd__nand3_1
Xhold919 top_inst.axis_out_inst.out_buff_data\[58\] VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16046_ _08532_ _08630_ _08629_ VGND VGND VPWR VPWR _08653_ sky130_fd_sc_hd__o21a_1
XFILLER_0_177_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13258_ _06032_ _06034_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__nor2_1
XFILLER_0_237_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12209_ top_inst.axis_out_inst.out_buff_data\[30\] _05129_ VGND VGND VPWR VPWR _05134_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_62_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13189_ _05959_ _05961_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19805_ _01600_ _01602_ _01630_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__a21o_1
X_17997_ _10499_ _10462_ VGND VGND VPWR VPWR _10500_ sky130_fd_sc_hd__nand2_1
XFILLER_0_236_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16948_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[10\] _09419_ VGND
+ VGND VPWR VPWR _09503_ sky130_fd_sc_hd__xnor2_1
X_19736_ _01563_ _01529_ VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__nor2_1
XFILLER_0_223_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16879_ _09427_ _09434_ _09435_ VGND VGND VPWR VPWR _09436_ sky130_fd_sc_hd__nand3_1
X_19667_ _01488_ _01495_ _01496_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__or3_4
XFILLER_0_126_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_232_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18618_ _10933_ _11056_ VGND VGND VPWR VPWR _11077_ sky130_fd_sc_hd__nor2_1
X_19598_ _01389_ _01429_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18549_ _11008_ _11009_ VGND VGND VPWR VPWR _11010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21560_ _02875_ _02895_ _03254_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20511_ _02292_ _02293_ _02286_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21491_ _03167_ _03183_ _03224_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_975 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23230_ net553 _04713_ _04724_ _04717_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20442_ _02188_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_209_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23161_ _04654_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20373_ _02157_ _02158_ _02159_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__and3_1
XFILLER_0_144_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22112_ top_inst.deskew_buff_inst.col_input\[101\] _05731_ _03802_ _03803_ VGND VGND
+ VPWR VPWR _03804_ sky130_fd_sc_hd__a22o_1
X_23092_ _04644_ net37 _04867_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22043_ _03723_ _03734_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23994_ clknet_leaf_82_clk _00527_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_242_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22945_ net643 _04548_ _04560_ _04551_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_242_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22876_ net784 _04517_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__or2_1
X_24615_ clknet_leaf_32_clk _01148_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dfxtp_4
X_21827_ _03509_ _03545_ _03542_ _03547_ _03541_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__a32o_1
XFILLER_0_214_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12560_ _05352_ _05374_ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24546_ clknet_leaf_103_clk _01079_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21758_ _03481_ _03482_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20709_ _02486_ _02454_ _02456_ _06404_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__a31oi_1
X_24477_ clknet_leaf_38_clk _01010_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_12491_ _04861_ _05309_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__nor2_2
XFILLER_0_124_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21689_ _03389_ _03416_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__xor2_2
XFILLER_0_151_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14230_ _06937_ _06940_ VGND VGND VPWR VPWR _06942_ sky130_fd_sc_hd__and2_1
X_23428_ _04863_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__buf_2
XFILLER_0_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14161_ _06872_ _06874_ VGND VGND VPWR VPWR _06875_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23359_ net43 _04792_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13112_ _05741_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[5\] VGND
+ VGND VPWR VPWR _05892_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14092_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[3\]\[2\]
+ _06806_ VGND VGND VPWR VPWR _06807_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13043_ top_inst.grid_inst.data_path_wires\[1\]\[2\] _05738_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _05825_ sky130_fd_sc_hd__nand4_1
X_17920_ _10423_ _10424_ VGND VGND VPWR VPWR _10425_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17851_ _10317_ _10356_ VGND VGND VPWR VPWR _10358_ sky130_fd_sc_hd__or2_1
XFILLER_0_218_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16802_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _09360_ sky130_fd_sc_hd__inv_2
X_17782_ _10252_ _10250_ VGND VGND VPWR VPWR _10290_ sky130_fd_sc_hd__or2b_1
XFILLER_0_205_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14994_ _07608_ _07606_ _07629_ _07627_ VGND VGND VPWR VPWR _07649_ sky130_fd_sc_hd__nand4_2
XFILLER_0_79_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19521_ _01352_ _01353_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__nor2_2
X_16733_ net1081 _09266_ _09291_ _09293_ _07708_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__o221a_1
X_13945_ _06662_ _06663_ _06664_ _06665_ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__a31o_1
XFILLER_0_205_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19452_ _01247_ _01260_ _01285_ _01286_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__o211a_1
X_16664_ _09226_ _09227_ _09222_ VGND VGND VPWR VPWR _09228_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_220_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13876_ _06609_ _06610_ _06615_ VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18403_ _10812_ _10810_ VGND VGND VPWR VPWR _10868_ sky130_fd_sc_hd__and2b_1
X_15615_ _08211_ _08214_ VGND VGND VPWR VPWR _08234_ sky130_fd_sc_hd__nand2_1
X_12827_ _05633_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__buf_6
X_19383_ _01186_ _01192_ _01191_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_887 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16595_ _09143_ _09144_ _09169_ _09141_ VGND VGND VPWR VPWR _09170_ sky130_fd_sc_hd__a211o_1
XFILLER_0_189_1032 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18334_ _10592_ _10602_ _10797_ _10798_ VGND VGND VPWR VPWR _10800_ sky130_fd_sc_hd__nand4_2
XFILLER_0_127_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15546_ _08150_ _07639_ _08170_ _08166_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__o211a_1
X_12758_ top_inst.axis_in_inst.inbuf_bus\[4\] _05267_ _05566_ VGND VGND VPWR VPWR
+ _05567_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_189_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18265_ _10727_ _10732_ VGND VGND VPWR VPWR _10733_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15477_ _08088_ _08090_ _08117_ VGND VGND VPWR VPWR _08118_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_126_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12689_ _05284_ _05301_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17216_ _09748_ _09763_ VGND VGND VPWR VPWR _09764_ sky130_fd_sc_hd__xor2_1
XFILLER_0_170_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14428_ _07121_ _07122_ _07104_ _07105_ VGND VGND VPWR VPWR _07124_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_163_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18196_ _10664_ _10665_ VGND VGND VPWR VPWR _10666_ sky130_fd_sc_hd__nand2_1
XFILLER_0_181_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17147_ _09696_ _09691_ VGND VGND VPWR VPWR _09697_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14359_ _07064_ VGND VGND VPWR VPWR _07065_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold705 _00059_ VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold716 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[4\] VGND VGND
+ VPWR VPWR net898 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold727 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[8\] VGND
+ VGND VPWR VPWR net909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 top_inst.axis_out_inst.out_buff_data\[59\] VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17078_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[12\] _09628_ _09629_
+ VGND VGND VPWR VPWR _09630_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_1060 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold749 _00167_ VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16029_ _08603_ _08606_ _08605_ VGND VGND VPWR VPWR _08637_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_23_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_1244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_240_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19719_ _01500_ _01523_ _01546_ _01547_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20991_ _02733_ _02736_ _02757_ _01984_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__a31o_1
XFILLER_0_237_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22730_ _04398_ _04400_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__and2_1
XFILLER_0_177_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22661_ _04334_ _04335_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__and2_1
XFILLER_0_211_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24400_ clknet_leaf_39_clk net765 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21612_ _03339_ _03342_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22592_ _04267_ _04269_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__xor2_1
XFILLER_0_63_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24331_ clknet_leaf_6_clk _00864_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21543_ _03190_ _03192_ _03231_ _03237_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24262_ clknet_leaf_110_clk _00795_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_21474_ _02891_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[3\] _02878_
+ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23213_ net595 _04713_ _04715_ _04704_ VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__o211a_1
X_20425_ _02208_ _02209_ _02164_ _02166_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__a211o_1
XFILLER_0_160_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24193_ clknet_leaf_117_clk _00726_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23144_ net632 _04671_ _04674_ _04675_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__o211a_1
X_20356_ _02141_ _02142_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__or2_1
XFILLER_0_219_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23075_ net17 _04628_ _04635_ _04632_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20287_ _01997_ _02007_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__nand2_2
XTAP_6226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22026_ _03720_ _03721_ _03715_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__a21o_1
XTAP_6259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold76 top_inst.axis_in_inst.inbuf_bus\[7\] VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold87 _00121_ VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11991_ _05009_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__clkbuf_2
Xhold98 top_inst.deskew_buff_inst.col_input\[49\] VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__dlygate4sd3_1
X_23977_ clknet_leaf_87_clk _00510_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13730_ _06433_ _06435_ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__or2_1
X_22928_ net991 _04548_ _04549_ _04551_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_211_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13661_ _06407_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__clkbuf_1
X_22859_ net809 _04504_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__or2_1
XFILLER_0_196_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15400_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[12\] _07924_ _07844_
+ VGND VGND VPWR VPWR _08043_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12612_ _05280_ _05297_ _05301_ _05273_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__a22oi_1
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16380_ _08669_ _08671_ _08697_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _08960_ sky130_fd_sc_hd__and4b_1
XFILLER_0_155_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13592_ _06327_ _06339_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15331_ _07970_ _07975_ VGND VGND VPWR VPWR _07976_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12543_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[0\]
+ _05286_ _05291_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__and4_1
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24529_ clknet_leaf_130_clk _01062_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_54_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18050_ _10548_ _10550_ VGND VGND VPWR VPWR _10551_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15262_ _07876_ _07882_ _07907_ VGND VGND VPWR VPWR _07908_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12474_ top_inst.skew_buff_inst.row\[0\].output_reg\[5\] top_inst.axis_in_inst.inbuf_bus\[5\]
+ net213 VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__mux2_4
XFILLER_0_152_956 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17001_ _09360_ _09377_ _09205_ _09209_ VGND VGND VPWR VPWR _09555_ sky130_fd_sc_hd__or4b_4
XFILLER_0_22_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14213_ top_inst.grid_inst.data_path_wires\[3\]\[4\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15193_ _07624_ _07622_ _07629_ _07627_ VGND VGND VPWR VPWR _07841_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 _10831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14144_ top_inst.grid_inst.data_path_wires\[3\]\[6\] top_inst.grid_inst.data_path_wires\[3\]\[5\]
+ _06648_ _06645_ VGND VGND VPWR VPWR _06858_ sky130_fd_sc_hd__and4_1
XFILLER_0_50_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14075_ _06751_ _06790_ VGND VGND VPWR VPWR _06791_ sky130_fd_sc_hd__xnor2_2
X_18952_ _11373_ _11374_ VGND VGND VPWR VPWR _11375_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13026_ _05803_ _05808_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__xnor2_1
X_17903_ _10407_ VGND VGND VPWR VPWR _10408_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18883_ _11300_ _11306_ VGND VGND VPWR VPWR _11307_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17834_ top_inst.grid_inst.data_path_wires\[11\]\[4\] _10056_ _10300_ top_inst.grid_inst.data_path_wires\[11\]\[3\]
+ VGND VGND VPWR VPWR _10341_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_59_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14977_ _07615_ _06647_ _07636_ _07618_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17765_ _10271_ _10273_ VGND VGND VPWR VPWR _10274_ sky130_fd_sc_hd__nand2_1
XFILLER_0_238_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer19 _09519_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19504_ _01287_ _01335_ _01337_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16716_ _09274_ _09275_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[4\]
+ VGND VGND VPWR VPWR _09277_ sky130_fd_sc_hd__a21oi_1
X_13928_ _06652_ _06641_ VGND VGND VPWR VPWR _06653_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17696_ _10032_ _10029_ _10052_ _10050_ VGND VGND VPWR VPWR _10206_ sky130_fd_sc_hd__nand4_2
XFILLER_0_77_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16647_ top_inst.skew_buff_inst.row\[2\].output_reg\[6\] top_inst.axis_in_inst.inbuf_bus\[22\]
+ _05266_ VGND VGND VPWR VPWR _09214_ sky130_fd_sc_hd__mux2_4
XFILLER_0_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19435_ _11697_ _11687_ _11692_ _11693_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13859_ _06555_ _06599_ VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_230_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16578_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[15\] _08975_ VGND
+ VGND VPWR VPWR _09153_ sky130_fd_sc_hd__xnor2_2
X_19366_ _11683_ net233 _11695_ _11678_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18317_ _10781_ _10782_ _05353_ VGND VGND VPWR VPWR _10784_ sky130_fd_sc_hd__a21o_1
X_15529_ _08137_ _07639_ _08158_ _08142_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__o211a_1
X_19297_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _11697_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18248_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[5\] _10693_ _10694_
+ VGND VGND VPWR VPWR _10716_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_154_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18179_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[3\] _10648_ _10649_
+ VGND VGND VPWR VPWR _10650_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold502 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[29\] VGND
+ VGND VPWR VPWR net684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold513 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[29\] VGND
+ VGND VPWR VPWR net695 sky130_fd_sc_hd__dlygate4sd3_1
X_20210_ _02009_ _11689_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold524 top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[31\] VGND VGND
+ VPWR VPWR net706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21190_ _02930_ _02931_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__or2_1
Xhold535 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[0\] VGND
+ VGND VPWR VPWR net717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[1\] VGND VGND
+ VPWR VPWR net728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold557 top_inst.axis_out_inst.out_buff_data\[119\] VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20141_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[30\] _01764_ VGND
+ VGND VPWR VPWR _01952_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold568 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[3\] VGND
+ VGND VPWR VPWR net750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[2\] VGND VGND
+ VPWR VPWR net761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_216_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20072_ top_inst.deskew_buff_inst.col_input\[26\] _05730_ VGND VGND VPWR VPWR _01887_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_141_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23900_ clknet_leaf_51_clk _00433_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_176_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1063 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23831_ clknet_leaf_93_clk _00364_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23762_ clknet_leaf_66_clk _00295_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_170_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20974_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[25\] _02468_ VGND
+ VGND VPWR VPWR _02742_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22713_ _04364_ _04382_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23693_ clknet_leaf_119_clk _00226_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22644_ _04317_ _04318_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22575_ _04210_ _04234_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24314_ clknet_leaf_1_clk _00847_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[89\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21526_ _02875_ _02893_ _03214_ _03258_ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__a31o_1
XFILLER_0_173_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24245_ clknet_leaf_126_clk _00778_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21457_ _03072_ _03112_ _03157_ _03191_ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__a31o_1
XFILLER_0_142_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12190_ net352 _05110_ _05122_ _05114_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__o211a_1
X_20408_ top_inst.grid_inst.data_path_wires\[16\]\[6\] _02009_ _02192_ _02193_ VGND
+ VGND VPWR VPWR _02194_ sky130_fd_sc_hd__nand4_2
X_24176_ clknet_leaf_27_clk _00709_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_21388_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[8\] _03122_ _03123_
+ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23127_ net422 _04656_ _04665_ _04662_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput44 net44 VGND VGND VPWR VPWR output_tdata[105] sky130_fd_sc_hd__clkbuf_4
XTAP_6001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20339_ _02125_ _02126_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__and2_2
XTAP_6012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput55 net55 VGND VGND VPWR VPWR output_tdata[115] sky130_fd_sc_hd__clkbuf_4
XTAP_6023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput66 net66 VGND VGND VPWR VPWR output_tdata[125] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_179_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput77 net77 VGND VGND VPWR VPWR output_tdata[1] sky130_fd_sc_hd__buf_2
Xoutput88 net88 VGND VGND VPWR VPWR output_tdata[2] sky130_fd_sc_hd__clkbuf_4
X_23058_ net9 _04615_ _04625_ _04619_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__o211a_1
XTAP_6045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput99 net99 VGND VGND VPWR VPWR output_tdata[3] sky130_fd_sc_hd__buf_2
XTAP_6067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14900_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[15\] _07364_ _07280_
+ VGND VGND VPWR VPWR _07583_ sky130_fd_sc_hd__a21oi_1
XTAP_5333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22009_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _03709_ sky130_fd_sc_hd__clkbuf_4
XTAP_6089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880_ _08484_ _08491_ VGND VGND VPWR VPWR _08492_ sky130_fd_sc_hd__nand2_1
XTAP_5355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14831_ _07484_ _07516_ VGND VGND VPWR VPWR _07517_ sky130_fd_sc_hd__xor2_2
XTAP_5388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[1\] _10064_ _10065_
+ VGND VGND VPWR VPWR _10066_ sky130_fd_sc_hd__nand3_1
X_14762_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[11\] _07364_ _07280_
+ VGND VGND VPWR VPWR _07449_ sky130_fd_sc_hd__a21o_1
XTAP_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ top_inst.axis_out_inst.out_buff_data\[57\] _04996_ VGND VGND VPWR VPWR _05000_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_99_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_230_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16501_ _09078_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13713_ top_inst.grid_inst.data_path_wires\[2\]\[7\] _06210_ _06208_ VGND VGND VPWR
+ VPWR _06458_ sky130_fd_sc_hd__and3_2
X_17481_ _09194_ _09189_ VGND VGND VPWR VPWR _10015_ sky130_fd_sc_hd__nand2_1
XTAP_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14693_ _07083_ _07082_ _07379_ _07380_ VGND VGND VPWR VPWR _07382_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16432_ _08676_ _08695_ VGND VGND VPWR VPWR _09011_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19220_ _11633_ _11634_ VGND VGND VPWR VPWR _11636_ sky130_fd_sc_hd__nand2_1
X_13644_ _06387_ _06388_ _06390_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_224_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19151_ _11557_ _11529_ _11568_ VGND VGND VPWR VPWR _11569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16363_ _08937_ _08943_ VGND VGND VPWR VPWR _08944_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ _05325_ _06323_ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__or2_1
XFILLER_0_171_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18102_ _10587_ _04859_ VGND VGND VPWR VPWR _10588_ sky130_fd_sc_hd__nand2_1
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_240_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15314_ _07957_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[7\] _07640_
+ top_inst.grid_inst.data_path_wires\[6\]\[5\] VGND VGND VPWR VPWR _07959_ sky130_fd_sc_hd__a22o_1
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12526_ _05321_ _05330_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19082_ _11460_ _11463_ _11501_ VGND VGND VPWR VPWR _11502_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_1143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16294_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _08876_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18033_ _10488_ _10510_ _10508_ VGND VGND VPWR VPWR _10535_ sky130_fd_sc_hd__o21a_1
X_15245_ _07887_ _07891_ VGND VGND VPWR VPWR _07892_ sky130_fd_sc_hd__xor2_2
X_12457_ top_inst.skew_buff_inst.row\[0\].output_reg\[2\] top_inst.axis_in_inst.inbuf_bus\[2\]
+ net213 VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__mux2_4
XFILLER_0_169_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15176_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _07824_ sky130_fd_sc_hd__inv_2
X_12388_ net807 _05230_ _05236_ _05234_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__o211a_1
XFILLER_0_238_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14127_ _06839_ _06841_ VGND VGND VPWR VPWR _06842_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19984_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[23\] _01764_ VGND
+ VGND VPWR VPWR _01802_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14058_ _06772_ _06773_ VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__xnor2_2
X_18935_ _11348_ _11357_ VGND VGND VPWR VPWR _11358_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_238_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13009_ _05777_ _05781_ _05792_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18866_ _11288_ _11289_ _11251_ _11250_ VGND VGND VPWR VPWR _11291_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_98_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1039 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17817_ _10279_ _10319_ _10323_ _10278_ VGND VGND VPWR VPWR _10324_ sky130_fd_sc_hd__a22o_1
XFILLER_0_222_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18797_ _11222_ _11223_ VGND VGND VPWR VPWR _11224_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17748_ _10254_ _10256_ VGND VGND VPWR VPWR _10257_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17679_ _10188_ _10189_ VGND VGND VPWR VPWR _10190_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19418_ _01250_ _01251_ _01253_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__nand3_1
X_20690_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[14\] _02468_ VGND
+ VGND VPWR VPWR _02469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19349_ _11683_ _11687_ _11692_ _11678_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22360_ _04013_ _04045_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21311_ _03047_ _03048_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__xor2_1
X_22291_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[9\] _03937_ _03938_
+ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_241_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24030_ clknet_leaf_41_clk _00563_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21242_ _02926_ _02947_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_206_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold310 top_inst.axis_out_inst.out_buff_data\[30\] VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 top_inst.deskew_buff_inst.col_input\[82\] VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[3\] VGND
+ VGND VPWR VPWR net514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 _00063_ VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold354 _00274_ VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__dlygate4sd3_1
X_21173_ _02914_ _02915_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__xor2_1
Xhold365 _00142_ VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[4\] VGND
+ VGND VPWR VPWR net558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold387 _00271_ VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__dlygate4sd3_1
X_20124_ _01563_ _01935_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__nor2_1
Xhold398 top_inst.valid_pipe\[0\] VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20055_ _01845_ _01848_ _01847_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23814_ clknet_leaf_72_clk _00347_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23745_ clknet_leaf_122_clk _00278_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20957_ _02528_ _02717_ _02724_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__nand3_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23676_ clknet_leaf_116_clk net427 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20888_ _02641_ _02659_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22627_ _04302_ _04303_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13360_ _06102_ _06101_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22558_ _04137_ _04223_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__nor2_1
XFILLER_0_187_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12311_ net916 _05191_ _05192_ _05182_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21509_ _03203_ _03202_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__or2b_1
XFILLER_0_224_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13291_ _06065_ _06066_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__nor2_1
X_22489_ _04143_ _04134_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1063 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15030_ _07668_ _07662_ _07680_ VGND VGND VPWR VPWR _07683_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12242_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[12\] _05143_
+ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__or2_1
X_24228_ clknet_leaf_112_clk _00761_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[16\]\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_210_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12173_ top_inst.axis_out_inst.out_buff_data\[15\] _05102_ VGND VGND VPWR VPWR _05113_
+ sky130_fd_sc_hd__or2_1
X_24159_ clknet_leaf_9_clk _00692_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16981_ _09534_ _09532_ VGND VGND VPWR VPWR _09536_ sky130_fd_sc_hd__and2b_1
XFILLER_0_236_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_1247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18720_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _11156_ sky130_fd_sc_hd__clkbuf_4
XTAP_5130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15932_ _08540_ _08542_ VGND VGND VPWR VPWR _08543_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_235_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15863_ _08475_ VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18651_ _11107_ _11108_ VGND VGND VPWR VPWR _11109_ sky130_fd_sc_hd__nand2_1
XTAP_5185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14814_ _07459_ _07499_ VGND VGND VPWR VPWR _07500_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_203_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ top_inst.grid_inst.data_path_wires\[11\]\[0\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[11\]\[1\]
+ VGND VGND VPWR VPWR _10115_ sky130_fd_sc_hd__a22o_1
XFILLER_0_235_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_204_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15794_ _08405_ _08407_ VGND VGND VPWR VPWR _08408_ sky130_fd_sc_hd__and2_1
X_18582_ _11041_ VGND VGND VPWR VPWR _11042_ sky130_fd_sc_hd__inv_2
XTAP_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14745_ _07431_ _07432_ VGND VGND VPWR VPWR _07433_ sky130_fd_sc_hd__nand2_1
XTAP_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ _10032_ _10046_ _10053_ _10049_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__o211a_1
XTAP_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ net864 _04977_ _04989_ _04981_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17464_ _09992_ _09985_ _09998_ _09999_ VGND VGND VPWR VPWR _10000_ sky130_fd_sc_hd__a211o_1
XFILLER_0_157_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14676_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[9\] _07364_ _07280_
+ VGND VGND VPWR VPWR _07365_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11888_ net886 _04938_ _04950_ _04942_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16415_ _08992_ _08994_ VGND VGND VPWR VPWR _08995_ sky130_fd_sc_hd__nand2_1
X_19203_ _11585_ _11615_ _11618_ VGND VGND VPWR VPWR _11619_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_117_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13627_ _06371_ _06373_ VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__xnor2_1
X_17395_ _09915_ _09916_ VGND VGND VPWR VPWR _09934_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_8__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_4_8__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_16346_ _08925_ _08926_ VGND VGND VPWR VPWR _08927_ sky130_fd_sc_hd__xor2_1
X_19134_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[13\] _11469_ VGND
+ VGND VPWR VPWR _11552_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13558_ top_inst.grid_inst.data_path_wires\[2\]\[5\] _06202_ _06200_ _06195_ VGND
+ VGND VPWR VPWR _06307_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_137_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12509_ _05326_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__clkbuf_16
X_19065_ _11482_ _11484_ VGND VGND VPWR VPWR _11485_ sky130_fd_sc_hd__nor2_1
X_16277_ _08857_ _08859_ VGND VGND VPWR VPWR _08860_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13489_ _06239_ _06240_ _05336_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15228_ _07825_ _07827_ _07823_ VGND VGND VPWR VPWR _07875_ sky130_fd_sc_hd__o21ba_1
X_18016_ _10071_ _10517_ _10518_ _10448_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15159_ _07805_ _07807_ VGND VGND VPWR VPWR _07808_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19967_ _01778_ _01785_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18918_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[8\] _11340_ VGND
+ VGND VPWR VPWR _11341_ sky130_fd_sc_hd__xnor2_1
X_19898_ _01562_ _01699_ _01719_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_207_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18849_ _11272_ _11273_ VGND VGND VPWR VPWR _11274_ sky130_fd_sc_hd__nor2_1
XFILLER_0_241_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21860_ _03578_ _03579_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20811_ _02556_ _02572_ _02585_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_222_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21791_ _03491_ _03494_ _03513_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_188_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23530_ clknet_leaf_140_clk net525 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20742_ _02518_ _02501_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23461_ net517 _04864_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20673_ net837 _01386_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22412_ _04060_ _04095_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__xor2_1
X_23392_ net59 _04805_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22343_ _04027_ _04028_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22274_ _03902_ _03910_ _03961_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24013_ clknet_leaf_48_clk _00546_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_143_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold140 _00286_ VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__dlygate4sd3_1
X_21225_ _02862_ _02893_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold151 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[22\] VGND
+ VGND VPWR VPWR net333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold162 _00202_ VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold173 top_inst.deskew_buff_inst.col_input\[4\] VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold184 _00190_ VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 top_inst.axis_out_inst.out_buff_data\[67\] VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__dlygate4sd3_1
X_21156_ _02899_ _02900_ _06178_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_106_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20107_ _01918_ _01919_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__and2_1
X_21087_ _02840_ _02847_ _02849_ VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__o21a_1
XFILLER_0_176_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_232_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20038_ _01844_ _01852_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__or2_1
XFILLER_0_226_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ _05635_ _05629_ _05666_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_77_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ net742 _04903_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__or2_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12791_ _05596_ _05598_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__nand2_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21989_ top_inst.grid_inst.data_path_wires\[18\]\[7\] VGND VGND VPWR VPWR _03695_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_150_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14530_ _07185_ _07222_ _07188_ _07161_ VGND VGND VPWR VPWR _07223_ sky130_fd_sc_hd__a2bb2o_2
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11742_ _04863_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__buf_2
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23728_ clknet_leaf_121_clk _00261_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_230_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _07154_ _07155_ VGND VGND VPWR VPWR _07156_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23659_ clknet_leaf_132_clk net527 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_230_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16200_ _08736_ _08758_ _08784_ VGND VGND VPWR VPWR _08785_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13412_ _05260_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__buf_2
XFILLER_0_37_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17180_ _09417_ _09418_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[16\]
+ VGND VGND VPWR VPWR _09729_ sky130_fd_sc_hd__or3b_1
XFILLER_0_92_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14392_ _05260_ VGND VGND VPWR VPWR _07092_ sky130_fd_sc_hd__buf_4
XFILLER_0_37_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16131_ _08717_ _08718_ VGND VGND VPWR VPWR _08719_ sky130_fd_sc_hd__and2_1
X_13343_ _05751_ _06082_ _06115_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__nor3_1
XFILLER_0_49_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16062_ _08137_ _08663_ _08665_ _08666_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13274_ _06048_ _06049_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15013_ _06848_ _07665_ _07666_ _07643_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12225_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[4\] _05143_
+ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19821_ _01627_ _01622_ _01645_ _10957_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__a31o_1
XFILLER_0_241_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12156_ top_inst.axis_out_inst.out_buff_data\[7\] _05102_ VGND VGND VPWR VPWR _05104_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_124_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19752_ _01577_ _01578_ _01579_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__nand3_1
X_16964_ _09516_ _09517_ _09509_ VGND VGND VPWR VPWR _09519_ sky130_fd_sc_hd__a21o_1
X_12087_ net520 _05063_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__or2_1
XFILLER_0_235_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18703_ _10589_ _11142_ _11144_ _11137_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__o211a_1
X_15915_ _08484_ _08524_ VGND VGND VPWR VPWR _08526_ sky130_fd_sc_hd__or2_1
XFILLER_0_223_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19683_ _01474_ _01470_ _01511_ _10957_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__a31o_1
X_16895_ _08870_ _09450_ _09451_ _09231_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18634_ _11075_ _11092_ VGND VGND VPWR VPWR _11093_ sky130_fd_sc_hd__xnor2_1
XTAP_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _08413_ _08411_ VGND VGND VPWR VPWR _08459_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18565_ _11024_ _11025_ VGND VGND VPWR VPWR _11026_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12989_ _05317_ _05775_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__nand2_1
XTAP_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15777_ _08350_ _08351_ _08390_ VGND VGND VPWR VPWR _08392_ sky130_fd_sc_hd__nand3_1
XTAP_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17516_ _10040_ _10033_ _10041_ _10024_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14728_ net1123 VGND VGND VPWR VPWR _07416_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18496_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[11\] _10364_ _10956_
+ _10958_ _09886_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14659_ _07346_ _07348_ VGND VGND VPWR VPWR _07349_ sky130_fd_sc_hd__xnor2_4
X_17447_ _09965_ _09983_ VGND VGND VPWR VPWR _09984_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17378_ _09917_ VGND VGND VPWR VPWR _09918_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19117_ _11511_ _11535_ VGND VGND VPWR VPWR _11536_ sky130_fd_sc_hd__or2b_1
X_16329_ _08857_ _08859_ VGND VGND VPWR VPWR _08911_ sky130_fd_sc_hd__and2b_1
XFILLER_0_125_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_207_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19048_ _11431_ _11434_ _11467_ VGND VGND VPWR VPWR _11468_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21010_ _02754_ _02776_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_214_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22961_ net734 _04562_ _04569_ _04564_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21912_ _03453_ _03617_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__or2b_1
XFILLER_0_74_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22892_ _06619_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__buf_2
XFILLER_0_218_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24631_ clknet_leaf_25_clk _01164_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[107\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21843_ _03550_ _03562_ _03552_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__or3_1
XFILLER_0_214_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24562_ clknet_leaf_137_clk _01095_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21774_ _03496_ _03497_ VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23513_ clknet_leaf_137_clk _00046_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20725_ _02461_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__clkbuf_4
X_24493_ clknet_leaf_125_clk _01026_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_92_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23444_ net627 _04840_ _04843_ _04844_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_1434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20656_ _02428_ _02435_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__xor2_1
XFILLER_0_191_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23375_ net51 _04805_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20587_ _02001_ _02018_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22326_ _03969_ _04004_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22257_ _03939_ _03944_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__xor2_2
XFILLER_0_225_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12010_ net871 _05018_ _05020_ _05008_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__o211a_1
X_21208_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[3\] _02928_ _02929_
+ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_218_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22188_ _03876_ _03877_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21139_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _02889_ sky130_fd_sc_hd__buf_2
XFILLER_0_206_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_217_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13961_ _06664_ _06679_ VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__or2_1
XFILLER_0_205_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12912_ _05715_ _05716_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__nand2_1
X_15700_ _08275_ _08315_ VGND VGND VPWR VPWR _08316_ sky130_fd_sc_hd__xor2_1
X_16680_ _09229_ _09242_ VGND VGND VPWR VPWR _09243_ sky130_fd_sc_hd__nand2_1
XFILLER_0_198_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13892_ _06188_ _06192_ _06627_ _06446_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__o211a_1
XFILLER_0_241_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12843_ _05608_ _05649_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__xnor2_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15631_ _08139_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[2\] _08227_
+ _08200_ _08164_ VGND VGND VPWR VPWR _08249_ sky130_fd_sc_hd__a32o_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18350_ _10760_ _10774_ _10815_ VGND VGND VPWR VPWR _10816_ sky130_fd_sc_hd__o21a_1
X_15562_ _05787_ VGND VGND VPWR VPWR _08183_ sky130_fd_sc_hd__buf_8
X_12774_ _05507_ _05581_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__nand2_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _07204_ _07205_ VGND VGND VPWR VPWR _07206_ sky130_fd_sc_hd__nor2_1
X_17301_ _09842_ _09843_ VGND VGND VPWR VPWR _09845_ sky130_fd_sc_hd__and2_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _08116_ _08118_ _08119_ _08132_ VGND VGND VPWR VPWR _08133_ sky130_fd_sc_hd__o31a_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18281_ _10641_ _10748_ VGND VGND VPWR VPWR _10749_ sky130_fd_sc_hd__and2_1
XFILLER_0_232_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17232_ _09759_ _09751_ VGND VGND VPWR VPWR _09779_ sky130_fd_sc_hd__or2b_1
X_14444_ _07136_ _07137_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[4\]
+ VGND VGND VPWR VPWR _07139_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_232_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17163_ _09699_ _09686_ _09711_ VGND VGND VPWR VPWR _09713_ sky130_fd_sc_hd__and3_1
XFILLER_0_181_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14375_ _07077_ VGND VGND VPWR VPWR _07078_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16114_ _08664_ _08683_ _08661_ _08686_ VGND VGND VPWR VPWR _08703_ sky130_fd_sc_hd__a22o_1
X_13326_ _06095_ _06100_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__xnor2_1
X_17094_ _09642_ _09643_ _09644_ VGND VGND VPWR VPWR _09646_ sky130_fd_sc_hd__a21o_1
Xhold909 top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[12\] VGND VGND
+ VPWR VPWR net1091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16045_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[15\] _08452_ _08373_
+ VGND VGND VPWR VPWR _08652_ sky130_fd_sc_hd__a21o_1
X_13257_ _05995_ _05997_ _06033_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12208_ net375 _05123_ _05133_ _05128_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__o211a_1
XFILLER_0_237_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13188_ _05966_ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19804_ _01562_ _01601_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12139_ top_inst.axis_out_inst.out_buff_data\[0\] _05089_ VGND VGND VPWR VPWR _05094_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_100_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_237_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17996_ _10040_ _10054_ VGND VGND VPWR VPWR _10499_ sky130_fd_sc_hd__and2_1
XFILLER_0_193_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19735_ _01562_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16947_ _09198_ _09219_ _09467_ _09466_ _09215_ VGND VGND VPWR VPWR _09502_ sky130_fd_sc_hd__a32o_1
XFILLER_0_223_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19666_ _01492_ _01493_ _01494_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__a21oi_1
X_16878_ _09431_ _09432_ _09433_ VGND VGND VPWR VPWR _09435_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18617_ _10969_ _11047_ _11049_ VGND VGND VPWR VPWR _11076_ sky130_fd_sc_hd__o21ai_1
X_15829_ _08399_ _08401_ _08398_ VGND VGND VPWR VPWR _08442_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_232_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19597_ _01390_ _01428_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_231_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18548_ _10969_ _11007_ VGND VGND VPWR VPWR _11009_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18479_ _10933_ _10941_ VGND VGND VPWR VPWR _10942_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20510_ _02286_ _02292_ _02293_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__nand3_1
XFILLER_0_145_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21490_ _03180_ _03182_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20441_ _02180_ _02182_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_1141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_892 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23160_ net830 _04671_ _04683_ _04675_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20372_ _02108_ _02116_ _02115_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_207_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22111_ _03777_ _03801_ _10831_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23091_ net33 VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22042_ _03070_ _03735_ _03736_ _03702_ VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23993_ clknet_leaf_79_clk _00526_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_242_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22944_ top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[1\] _04557_ VGND
+ VGND VPWR VPWR _04560_ sky130_fd_sc_hd__or2_1
XFILLER_0_223_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22875_ net707 _04509_ _04520_ _04511_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24614_ clknet_leaf_21_clk _01147_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_211_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21826_ _03519_ _03523_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_214_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24545_ clknet_leaf_100_clk _01078_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_144_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_144_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21757_ _03456_ _03480_ _03471_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__nand3_1
XFILLER_0_4_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20708_ _02454_ _02456_ _02486_ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__a21o_1
X_24476_ clknet_leaf_39_clk _01009_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_12490_ _05267_ _04856_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__or2_4
XFILLER_0_19_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21688_ _03414_ _03415_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__or2b_1
XFILLER_0_80_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23427_ net302 _04827_ _04834_ _04831_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20639_ _02389_ _02419_ VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__xor2_1
XFILLER_0_149_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_1098 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire169 _05879_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_46_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14160_ _06823_ _06832_ _06873_ VGND VGND VPWR VPWR _06874_ sky130_fd_sc_hd__a21oi_1
X_23358_ net872 _04791_ _04797_ _04795_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13111_ _05889_ _05890_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22309_ _03956_ _03958_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__nand2_1
X_14091_ top_inst.grid_inst.data_path_wires\[3\]\[1\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__and2b_1
X_23289_ net645 _04752_ _04758_ _04756_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13042_ top_inst.grid_inst.data_path_wires\[1\]\[1\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[1\]\[2\]
+ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__a22o_1
XFILLER_0_219_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17850_ _10317_ _10356_ VGND VGND VPWR VPWR _10357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_219_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16801_ _09359_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17781_ _10284_ _10288_ VGND VGND VPWR VPWR _10289_ sky130_fd_sc_hd__xor2_1
X_14993_ _07606_ _07629_ _07627_ _07608_ VGND VGND VPWR VPWR _07648_ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19520_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[0\]
+ _11707_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__and3_2
XFILLER_0_79_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16732_ _09289_ _09290_ _09292_ VGND VGND VPWR VPWR _09293_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13944_ _06643_ _06618_ VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19451_ _01283_ _01284_ net218 _01236_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_92_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16663_ _09224_ _09225_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[1\]
+ VGND VGND VPWR VPWR _09227_ sky130_fd_sc_hd__a21oi_1
X_13875_ _06611_ _06614_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_199_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18402_ _10846_ _10866_ VGND VGND VPWR VPWR _10867_ sky130_fd_sc_hd__xnor2_1
X_12826_ _05325_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__buf_8
X_15614_ _08230_ _08232_ VGND VGND VPWR VPWR _08233_ sky130_fd_sc_hd__xor2_2
XFILLER_0_202_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19382_ _01210_ _01211_ _01217_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__a21oi_2
X_16594_ _09165_ _09167_ VGND VGND VPWR VPWR _09169_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_1408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_202_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18333_ _10592_ _10602_ _10797_ _10798_ VGND VGND VPWR VPWR _10799_ sky130_fd_sc_hd__a22o_1
X_12757_ _05267_ top_inst.skew_buff_inst.row\[0\].output_reg\[4\] VGND VGND VPWR VPWR
+ _05566_ sky130_fd_sc_hd__and2b_1
XFILLER_0_189_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15545_ _08169_ _07641_ VGND VGND VPWR VPWR _08170_ sky130_fd_sc_hd__or2_1
XFILLER_0_173_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_135_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_135_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15476_ _08114_ _08115_ VGND VGND VPWR VPWR _08117_ sky130_fd_sc_hd__and2_1
X_18264_ _10730_ _10731_ VGND VGND VPWR VPWR _10732_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12688_ _05497_ _05498_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17215_ _09761_ _09762_ VGND VGND VPWR VPWR _09763_ sky130_fd_sc_hd__or2_1
X_14427_ _07104_ _07105_ _07121_ _07122_ VGND VGND VPWR VPWR _07123_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_115_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18195_ _10606_ _10585_ _10600_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _10665_ sky130_fd_sc_hd__nand4_1
XFILLER_0_71_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14358_ top_inst.skew_buff_inst.row\[1\].output_reg\[1\] top_inst.axis_in_inst.inbuf_bus\[9\]
+ net208 VGND VGND VPWR VPWR _07064_ sky130_fd_sc_hd__mux2_4
XFILLER_0_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17146_ _09665_ _09689_ VGND VGND VPWR VPWR _09696_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold706 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[2\] VGND
+ VGND VPWR VPWR net888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 _00906_ VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ _05748_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[7\] _05770_
+ _05750_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__and4b_1
XFILLER_0_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold728 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[26\] VGND
+ VGND VPWR VPWR net910 sky130_fd_sc_hd__dlygate4sd3_1
X_17077_ _09417_ VGND VGND VPWR VPWR _09629_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_204_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14289_ _06963_ _06632_ _06997_ VGND VGND VPWR VPWR _06999_ sky130_fd_sc_hd__nor3_1
Xhold739 top_inst.deskew_buff_inst.col_input\[69\] VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1072 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16028_ _08627_ _08635_ VGND VGND VPWR VPWR _08636_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1004 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_236_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17979_ _10449_ _10443_ _10482_ VGND VGND VPWR VPWR _10483_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_237_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19718_ _01544_ _01545_ _01531_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_240_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20990_ _02733_ _02736_ _02757_ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_1319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19649_ _11688_ _11709_ _01442_ _01441_ _11697_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22660_ _04315_ _04333_ _04328_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__nand3_1
XFILLER_0_133_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21611_ _03275_ _03340_ _03341_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22591_ _04268_ _04245_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_126_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_126_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24330_ clknet_leaf_7_clk _00863_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21542_ _03070_ _03273_ _03274_ _02909_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24261_ clknet_leaf_110_clk _00794_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21473_ _03205_ _03206_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23212_ net100 _04714_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__or2_1
X_20424_ _02164_ _02166_ _02208_ _02209_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__o211ai_2
X_24192_ clknet_leaf_47_clk _00725_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23143_ _04550_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20355_ _02102_ _02139_ _02140_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__nor3_1
XFILLER_0_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23074_ top_inst.axis_in_inst.inbuf_bus\[24\] _04629_ VGND VGND VPWR VPWR _04635_
+ sky130_fd_sc_hd__or2_1
XTAP_6216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20286_ net497 _05634_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22025_ _03718_ _03719_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[1\]
+ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__a21o_1
XTAP_6249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold77 _00981_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11990_ _04863_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__clkbuf_4
Xhold88 top_inst.deskew_buff_inst.col_input\[48\] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dlygate4sd3_1
X_23976_ clknet_leaf_87_clk _00509_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_242_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold99 _00120_ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22927_ _04550_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__buf_2
XFILLER_0_151_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13660_ _06364_ _06406_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22858_ net1034 _04509_ _04510_ _04511_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12611_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[0\]
+ _05296_ _05300_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__and4_1
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21809_ _03278_ _03530_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__nor2_1
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_117_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13591_ _06333_ _06338_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__xnor2_1
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22789_ _04420_ _04421_ _04441_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15330_ _07971_ _07974_ VGND VGND VPWR VPWR _07975_ sky130_fd_sc_hd__xor2_2
X_12542_ _05355_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__inv_2
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24528_ clknet_leaf_130_clk _01061_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15261_ _07875_ _07874_ VGND VGND VPWR VPWR _07907_ sky130_fd_sc_hd__or2b_1
XFILLER_0_4_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24459_ clknet_leaf_54_clk _00992_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_12473_ _05290_ _05292_ _05295_ _05261_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17000_ _09211_ _09214_ VGND VGND VPWR VPWR _09554_ sky130_fd_sc_hd__and2_1
X_14212_ _06924_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15192_ _07837_ _07839_ VGND VGND VPWR VPWR _07840_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_8 clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14143_ _06630_ _06648_ _06645_ _06632_ VGND VGND VPWR VPWR _06857_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_22_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14074_ _06783_ _06789_ VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__xnor2_2
X_18951_ _11370_ _11372_ VGND VGND VPWR VPWR _11374_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13025_ _05806_ _05807_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__nor2_1
X_17902_ _10368_ _10373_ _10371_ VGND VGND VPWR VPWR _10407_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18882_ _11301_ _11305_ VGND VGND VPWR VPWR _11306_ sky130_fd_sc_hd__xor2_1
XFILLER_0_123_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17833_ top_inst.grid_inst.data_path_wires\[11\]\[3\] _10059_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[6\]
+ top_inst.grid_inst.data_path_wires\[11\]\[4\] VGND VGND VPWR VPWR _10340_ sky130_fd_sc_hd__and4b_1
XTAP_6783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17764_ _10224_ _10225_ _10272_ VGND VGND VPWR VPWR _10273_ sky130_fd_sc_hd__a21o_1
XFILLER_0_221_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14976_ _07635_ _07075_ VGND VGND VPWR VPWR _07636_ sky130_fd_sc_hd__or2_1
XFILLER_0_234_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19503_ _01336_ _01334_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16715_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[4\] _09274_ _09275_
+ VGND VGND VPWR VPWR _09276_ sky130_fd_sc_hd__and3_1
X_13927_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _06652_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_221_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17695_ top_inst.grid_inst.data_path_wires\[11\]\[3\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[11\]\[4\]
+ VGND VGND VPWR VPWR _10205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19434_ _01266_ _01267_ _01261_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__a21o_1
X_16646_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _09213_ sky130_fd_sc_hd__buf_2
XFILLER_0_134_1352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13858_ _06597_ _06598_ VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12809_ _05507_ _05615_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19365_ _06168_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__buf_4
X_16577_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[14\] _08975_ _08896_
+ VGND VGND VPWR VPWR _09152_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_108_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_146_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13789_ _06486_ _06489_ _06487_ VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_128_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18316_ _10781_ _10782_ VGND VGND VPWR VPWR _10783_ sky130_fd_sc_hd__nor2_1
XFILLER_0_210_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15528_ _08157_ _07641_ VGND VGND VPWR VPWR _08158_ sky130_fd_sc_hd__or2_1
X_19296_ _11695_ VGND VGND VPWR VPWR _11696_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18247_ _10690_ _10698_ VGND VGND VPWR VPWR _10715_ sky130_fd_sc_hd__and2_1
XFILLER_0_182_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15459_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[15\] _07576_ VGND
+ VGND VPWR VPWR _08100_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18178_ _10585_ _10581_ _10600_ _10597_ VGND VGND VPWR VPWR _10649_ sky130_fd_sc_hd__nand4_1
XFILLER_0_25_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold503 _00036_ VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1000 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17129_ _09671_ _09679_ VGND VGND VPWR VPWR _09680_ sky130_fd_sc_hd__xor2_1
Xhold514 top_inst.deskew_buff_inst.col_input\[56\] VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[3\] VGND VGND
+ VPWR VPWR net707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold536 top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[4\] VGND VGND
+ VPWR VPWR net718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold547 top_inst.axis_out_inst.out_buff_data\[120\] VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__dlygate4sd3_1
X_20140_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[29\] _01761_ _01762_
+ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__a21o_1
Xhold558 top_inst.deskew_buff_inst.col_input\[114\] VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold569 top_inst.axis_out_inst.out_buff_data\[125\] VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20071_ _01884_ _01864_ _01867_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__or3_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23830_ clknet_leaf_94_clk _00363_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_225_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23761_ clknet_leaf_122_clk net301 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20973_ _02643_ _02723_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__nand2_1
XFILLER_0_240_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22712_ _09787_ _04383_ _04384_ _03929_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23692_ clknet_leaf_120_clk _00225_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22643_ _04317_ _04318_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_857 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22574_ _04251_ _04252_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24313_ clknet_leaf_1_clk _00846_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[88\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21525_ _02873_ _02895_ _03212_ VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24244_ clknet_leaf_125_clk _00777_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_21456_ _03117_ _03115_ _03156_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_224_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20407_ top_inst.grid_inst.data_path_wires\[16\]\[5\] top_inst.grid_inst.data_path_wires\[16\]\[4\]
+ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[3\] _02051_ VGND VGND
+ VPWR VPWR _02193_ sky130_fd_sc_hd__nand4_4
XFILLER_0_189_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24175_ clknet_leaf_27_clk _00708_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21387_ _03077_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__clkbuf_4
X_23126_ net110 _04659_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__or2_1
X_20338_ _02100_ _02101_ _02124_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__nand3_1
XTAP_6002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput45 net45 VGND VGND VPWR VPWR output_tdata[106] sky130_fd_sc_hd__buf_2
XTAP_6013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput56 net56 VGND VGND VPWR VPWR output_tdata[116] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput67 net67 VGND VGND VPWR VPWR output_tdata[126] sky130_fd_sc_hd__clkbuf_4
XTAP_6024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput78 net78 VGND VGND VPWR VPWR output_tdata[20] sky130_fd_sc_hd__clkbuf_4
X_23057_ net991 _04616_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__or2_1
XTAP_6035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20269_ _01995_ _02007_ _02056_ _02058_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__nand4_2
XTAP_5312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput89 net89 VGND VGND VPWR VPWR output_tdata[30] sky130_fd_sc_hd__buf_2
XTAP_6057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22008_ _03688_ _05270_ _03708_ _03702_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__o211a_1
XTAP_6079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14830_ _07514_ _07515_ VGND VGND VPWR VPWR _07516_ sky130_fd_sc_hd__nand2_1
XTAP_5378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14761_ _07405_ _07408_ _07447_ VGND VGND VPWR VPWR _07448_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_192_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11973_ net814 _04990_ _04999_ _04995_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__o211a_1
XTAP_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23959_ clknet_leaf_89_clk _00492_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16500_ _08831_ _09077_ VGND VGND VPWR VPWR _09078_ sky130_fd_sc_hd__and2_1
XTAP_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _06455_ _06456_ VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__xor2_1
X_14692_ _07083_ _07082_ _07379_ _07380_ VGND VGND VPWR VPWR _07381_ sky130_fd_sc_hd__nand4_1
X_17480_ _09990_ _10000_ _10008_ VGND VGND VPWR VPWR _10014_ sky130_fd_sc_hd__and3_1
XFILLER_0_169_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16431_ _09008_ _09009_ VGND VGND VPWR VPWR _09010_ sky130_fd_sc_hd__and2b_1
XFILLER_0_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13643_ _06384_ _06345_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19150_ _11566_ _11567_ VGND VGND VPWR VPWR _11568_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16362_ _08938_ _08942_ VGND VGND VPWR VPWR _08943_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13574_ _06320_ _06321_ _06289_ _06285_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__o211a_1
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18101_ top_inst.grid_inst.data_path_wires\[12\]\[4\] VGND VGND VPWR VPWR _10587_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12525_ _05273_ _05287_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__nand2_1
X_15313_ top_inst.grid_inst.data_path_wires\[6\]\[5\] _07957_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[7\]
+ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[6\] VGND VGND VPWR VPWR
+ _07958_ sky130_fd_sc_hd__and4_1
XFILLER_0_109_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16293_ top_inst.grid_inst.data_path_wires\[8\]\[1\] top_inst.grid_inst.data_path_wires\[8\]\[2\]
+ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _08875_ sky130_fd_sc_hd__and4b_1
XFILLER_0_147_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19081_ _11457_ _11500_ VGND VGND VPWR VPWR _11501_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_240_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18032_ _10522_ _10533_ VGND VGND VPWR VPWR _10534_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12456_ _05270_ _05279_ _05281_ _05261_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__o211a_1
X_15244_ _07889_ _07890_ VGND VGND VPWR VPWR _07891_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15175_ top_inst.grid_inst.data_path_wires\[6\]\[1\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[7\]
+ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[6\]\[2\]
+ VGND VGND VPWR VPWR _07823_ sky130_fd_sc_hd__and4b_1
XFILLER_0_23_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12387_ net357 _05235_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14126_ _06792_ _06794_ _06840_ VGND VGND VPWR VPWR _06841_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_123_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_205_1364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19983_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[22\] _01761_ _01762_
+ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__a21o_1
XFILLER_0_238_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14057_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[5\] _06624_ VGND
+ VGND VPWR VPWR _06773_ sky130_fd_sc_hd__nand2_1
X_18934_ _11354_ _11356_ VGND VGND VPWR VPWR _11357_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13008_ top_inst.grid_inst.data_path_wires\[1\]\[3\] top_inst.grid_inst.data_path_wires\[1\]\[2\]
+ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__and4_1
X_18865_ _11251_ _11250_ _11288_ _11289_ VGND VGND VPWR VPWR _11290_ sky130_fd_sc_hd__and4bb_1
XTAP_6580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17816_ _10271_ _10273_ _10319_ VGND VGND VPWR VPWR _10323_ sky130_fd_sc_hd__a21o_1
XFILLER_0_206_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18796_ _11197_ _11198_ _11200_ _11201_ _11194_ VGND VGND VPWR VPWR _11223_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17747_ _10209_ _10215_ _10255_ VGND VGND VPWR VPWR _10256_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_234_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14959_ top_inst.grid_inst.data_path_wires\[6\]\[7\] VGND VGND VPWR VPWR _07624_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_221_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17678_ _10099_ _10121_ _10146_ _10150_ VGND VGND VPWR VPWR _10189_ sky130_fd_sc_hd__o31a_1
XFILLER_0_203_983 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19417_ _01195_ _01222_ _01252_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16629_ _09198_ _09199_ VGND VGND VPWR VPWR _09200_ sky130_fd_sc_hd__or2_1
XFILLER_0_174_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19348_ _01184_ _01185_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_1057 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19279_ net190 VGND VGND VPWR VPWR _11682_ sky130_fd_sc_hd__buf_2
XFILLER_0_150_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21310_ _02873_ _02887_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22290_ _03940_ _03941_ _03942_ _03944_ _03939_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__a32o_1
XFILLER_0_131_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_562 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold300 _00073_ VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__dlygate4sd3_1
X_21241_ _02964_ _02980_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__xor2_2
Xhold311 top_inst.axis_out_inst.out_buff_data\[32\] VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold322 _00057_ VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold333 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[14\] VGND
+ VGND VPWR VPWR net515 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold344 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[25\] VGND
+ VGND VPWR VPWR net526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 top_inst.axis_out_inst.out_buff_data\[82\] VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__dlygate4sd3_1
X_21172_ _02903_ _02904_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__nand2_1
XFILLER_0_229_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold366 top_inst.axis_out_inst.out_buff_data\[25\] VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 top_inst.deskew_buff_inst.col_input\[62\] VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__buf_1
X_20123_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[29\] _01764_ VGND
+ VGND VPWR VPWR _01935_ sky130_fd_sc_hd__xnor2_1
Xhold388 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[14\] VGND
+ VGND VPWR VPWR net570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 top_inst.deskew_buff_inst.col_input\[97\] VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__buf_1
XFILLER_0_110_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20054_ _01831_ _01868_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23813_ clknet_leaf_72_clk _00346_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23744_ clknet_leaf_127_clk net516 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20956_ _02528_ _02717_ _02724_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__a21o_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23675_ clknet_leaf_116_clk net465 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20887_ _02629_ _02658_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__xnor2_1
X_22626_ _04284_ _04301_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22557_ net923 _03528_ _04235_ _04236_ _09806_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__o221a_1
XFILLER_0_63_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12310_ net572 _05183_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21508_ _03226_ _03200_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__or2b_1
XFILLER_0_84_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13290_ _05945_ _06064_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__and2_1
X_22488_ _04162_ _04169_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12241_ net420 _05151_ _05152_ _05141_ VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__o211a_1
X_24227_ clknet_leaf_113_clk _00760_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[16\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21439_ top_inst.grid_inst.data_path_wires\[17\]\[4\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1097 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24158_ clknet_leaf_9_clk _00691_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12172_ net692 _05110_ _05112_ _05101_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__o211a_1
X_23109_ top_inst.axis_out_inst.out_buff_enabled _05323_ VGND VGND VPWR VPWR _04653_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_219_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16980_ _09532_ _09534_ VGND VGND VPWR VPWR _09535_ sky130_fd_sc_hd__or2b_1
XFILLER_0_21_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24089_ clknet_leaf_97_clk _00622_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15931_ _08498_ _08501_ _08541_ VGND VGND VPWR VPWR _08542_ sky130_fd_sc_hd__a21bo_1
XTAP_5131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18650_ _11079_ _11082_ _11106_ VGND VGND VPWR VPWR _11108_ sky130_fd_sc_hd__or3_1
XTAP_5175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15862_ _08197_ _08474_ VGND VGND VPWR VPWR _08475_ sky130_fd_sc_hd__and2_1
XTAP_5186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17601_ _10027_ _10047_ VGND VGND VPWR VPWR _10114_ sky130_fd_sc_hd__nand2_1
X_14813_ _07497_ _07498_ VGND VGND VPWR VPWR _07499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_204_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18581_ _11006_ _11010_ _11008_ VGND VGND VPWR VPWR _11041_ sky130_fd_sc_hd__a21o_1
XFILLER_0_235_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ _08406_ VGND VGND VPWR VPWR _08407_ sky130_fd_sc_hd__inv_2
XFILLER_0_192_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17532_ _10052_ _09199_ VGND VGND VPWR VPWR _10053_ sky130_fd_sc_hd__or2_1
X_14744_ _07428_ _07429_ _07430_ VGND VGND VPWR VPWR _07432_ sky130_fd_sc_hd__a21o_1
XTAP_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ net796 _04982_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__or2_1
XTAP_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17463_ _09978_ _09997_ _09993_ VGND VGND VPWR VPWR _09999_ sky130_fd_sc_hd__nor3_1
XFILLER_0_50_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14675_ _07281_ VGND VGND VPWR VPWR _07364_ sky130_fd_sc_hd__clkbuf_4
X_11887_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[20\] _04943_
+ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19202_ _11578_ _11614_ VGND VGND VPWR VPWR _11618_ sky130_fd_sc_hd__or2b_1
X_16414_ _08872_ _08916_ _08955_ _08993_ VGND VGND VPWR VPWR _08994_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13626_ _06328_ _06329_ _06372_ VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_32_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17394_ _09922_ _09924_ VGND VGND VPWR VPWR _09933_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19133_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[12\] _11469_ _11387_
+ VGND VGND VPWR VPWR _11551_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16345_ _08877_ _08879_ _08875_ VGND VGND VPWR VPWR _08926_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_109_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13557_ _06195_ top_inst.grid_inst.data_path_wires\[2\]\[5\] _06202_ _06200_ VGND
+ VGND VPWR VPWR _06306_ sky130_fd_sc_hd__and4_1
XFILLER_0_171_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19064_ _11145_ _11161_ _11480_ _11483_ VGND VGND VPWR VPWR _11484_ sky130_fd_sc_hd__o2bb2a_1
X_12508_ _05325_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__buf_8
X_16276_ _08808_ _08812_ _08858_ VGND VGND VPWR VPWR _08859_ sky130_fd_sc_hd__o21ai_1
X_13488_ _06227_ _06238_ _06237_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__o21a_1
XFILLER_0_70_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18015_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[14\] _09494_ VGND
+ VGND VPWR VPWR _10518_ sky130_fd_sc_hd__or2_1
X_12439_ net186 VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__buf_6
X_15227_ _07872_ _07873_ VGND VGND VPWR VPWR _07874_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15158_ _07760_ _07806_ VGND VGND VPWR VPWR _07807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14109_ _06632_ _06785_ VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19966_ _01782_ _01784_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__xor2_2
X_15089_ _07739_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18917_ _11338_ _11339_ VGND VGND VPWR VPWR _11340_ sky130_fd_sc_hd__nor2_4
X_19897_ _01698_ _01700_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__or2b_1
XFILLER_0_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18848_ _11164_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[5\] top_inst.grid_inst.data_path_wires\[13\]\[1\]
+ top_inst.grid_inst.data_path_wires\[13\]\[0\] VGND VGND VPWR VPWR _11273_ sky130_fd_sc_hd__and4_1
XFILLER_0_101_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18779_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[3\] _05730_ VGND
+ VGND VPWR VPWR _11207_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20810_ _02583_ _02584_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_210_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21790_ _03279_ _03492_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20741_ _02462_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_212_1154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23460_ net260 _04859_ _04852_ _04844_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20672_ _02423_ _02451_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__xor2_1
XFILLER_0_174_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22411_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[13\] _03894_ VGND
+ VGND VPWR VPWR _04095_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23391_ net517 _04804_ _04815_ _04808_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_clk clknet_4_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_668 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22342_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[18\]\[5\]
+ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22273_ _03907_ _03909_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24012_ clknet_leaf_47_clk _00545_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_130_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21224_ _02950_ _02954_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__and2b_1
Xhold130 _00215_ VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold141 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[15\] VGND
+ VGND VPWR VPWR net323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 _00285_ VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[18\] VGND
+ VGND VPWR VPWR net345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 _00203_ VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold185 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[9\] VGND
+ VGND VPWR VPWR net367 sky130_fd_sc_hd__dlygate4sd3_1
X_21155_ _02862_ _02883_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_217_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold196 top_inst.axis_out_inst.out_buff_data\[36\] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_244_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20106_ _01563_ _01917_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_217_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21086_ _02827_ _02848_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__nor2_1
XFILLER_0_244_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_233_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_97_clk clknet_4_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_226_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20037_ _01844_ _01852_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__nand2_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ net522 _04898_ _04906_ _04902_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__o211a_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12790_ _05447_ _05449_ _05292_ _05597_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__or4_1
XFILLER_0_115_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21988_ _02875_ _02877_ _03694_ _03660_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11741_ _04862_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__buf_8
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20939_ _02681_ _02703_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__or2b_1
X_23727_ clknet_leaf_121_clk _00260_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14460_ net1125 _07152_ _07153_ VGND VGND VPWR VPWR _07155_ sky130_fd_sc_hd__o21bai_2
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23658_ clknet_leaf_135_clk _00191_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13411_ _06181_ _05262_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__or2_1
X_14391_ _05269_ _07090_ VGND VGND VPWR VPWR _07091_ sky130_fd_sc_hd__or2_1
X_22609_ _04245_ _04285_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23589_ clknet_4_8__leaf_clk _00122_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_clk clknet_4_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13342_ _05751_ _06082_ _06115_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__o21a_1
X_16130_ _08710_ _08716_ VGND VGND VPWR VPWR _08718_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13273_ _06009_ _06012_ _06010_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__o21ba_1
X_16061_ _07617_ VGND VGND VPWR VPWR _08666_ sky130_fd_sc_hd__buf_2
XFILLER_0_49_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15012_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[2\] _06168_ VGND
+ VGND VPWR VPWR _07666_ sky130_fd_sc_hd__or2_1
X_12224_ _05142_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_103_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19820_ _01627_ _01622_ _01645_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12155_ net402 _05097_ _05103_ _05101_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19751_ _01488_ _01540_ _01539_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__o21bai_1
X_16963_ _09509_ _09516_ net226 VGND VGND VPWR VPWR _09518_ sky130_fd_sc_hd__nand3_1
X_12086_ net445 _05058_ _05064_ _05062_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_88_clk clknet_4_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_198_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18702_ _11143_ _11133_ VGND VGND VPWR VPWR _11144_ sky130_fd_sc_hd__or2_1
X_15914_ _08484_ _08524_ VGND VGND VPWR VPWR _08525_ sky130_fd_sc_hd__nand2_1
X_19682_ _01474_ _01470_ _01511_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16894_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[8\] _07866_ VGND
+ VGND VPWR VPWR _09451_ sky130_fd_sc_hd__or2_1
XFILLER_0_204_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18633_ _11090_ _11091_ VGND VGND VPWR VPWR _11092_ sky130_fd_sc_hd__and2_1
XTAP_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ _08451_ _08457_ VGND VGND VPWR VPWR _08458_ sky130_fd_sc_hd__xnor2_1
XTAP_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18564_ _11012_ _10984_ _11023_ VGND VGND VPWR VPWR _11025_ sky130_fd_sc_hd__nand3_1
XTAP_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ _08350_ _08351_ _08390_ VGND VGND VPWR VPWR _08391_ sky130_fd_sc_hd__a21o_1
XFILLER_0_231_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12988_ _05734_ _05757_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__nand2_1
XTAP_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17515_ _10030_ _09219_ VGND VGND VPWR VPWR _10041_ sky130_fd_sc_hd__or2_1
XTAP_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14727_ _07328_ _07414_ VGND VGND VPWR VPWR _07415_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_169_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11939_ net999 _04977_ _04979_ _04968_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18495_ _10914_ _10917_ _10955_ _10957_ VGND VGND VPWR VPWR _10958_ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17446_ _09980_ _09982_ VGND VGND VPWR VPWR _09983_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14658_ _07299_ _07300_ _07347_ VGND VGND VPWR VPWR _07348_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_74_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13609_ _06293_ _06356_ _06315_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__a21oi_1
X_17377_ _09915_ _09916_ VGND VGND VPWR VPWR _09917_ sky130_fd_sc_hd__xor2_1
XFILLER_0_172_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_972 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14589_ _07279_ VGND VGND VPWR VPWR _07280_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_clk clknet_4_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_16
X_19116_ _11519_ _11534_ VGND VGND VPWR VPWR _11535_ sky130_fd_sc_hd__xor2_1
X_16328_ _08908_ _08909_ VGND VGND VPWR VPWR _08910_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19047_ _11433_ _11432_ VGND VGND VPWR VPWR _11467_ sky130_fd_sc_hd__or2b_1
XFILLER_0_140_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16259_ _08673_ _08688_ _08839_ _08840_ VGND VGND VPWR VPWR _08842_ sky130_fd_sc_hd__nand4_2
XFILLER_0_28_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_239_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19949_ _01763_ _01768_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__xor2_2
Xclkbuf_leaf_79_clk clknet_4_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22960_ top_inst.skew_buff_inst.row\[1\].output_reg\[0\] _04557_ VGND VGND VPWR VPWR
+ _04569_ sky130_fd_sc_hd__or2_1
XFILLER_0_241_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21911_ _03596_ _03616_ _03614_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__o21a_1
XFILLER_0_218_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22891_ net761 _04522_ _04529_ _04524_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24630_ clknet_leaf_25_clk _01163_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[106\]
+ sky130_fd_sc_hd__dfxtp_1
X_21842_ _03550_ _03552_ _03562_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_223_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24561_ clknet_leaf_137_clk _01094_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dfxtp_4
X_21773_ _03375_ _03478_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__nor2_1
XFILLER_0_210_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23512_ clknet_leaf_137_clk _00045_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_20724_ _02463_ _02501_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24492_ clknet_leaf_109_clk _01025_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_110_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23443_ _04869_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20655_ _02429_ _02434_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23374_ net423 _04804_ _04806_ _04795_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__o211a_1
X_20586_ _01999_ _02227_ _02367_ _02186_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__a22o_1
XFILLER_0_225_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22325_ _04011_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22256_ _03940_ _03943_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21207_ _02926_ _02947_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__xor2_2
XFILLER_0_197_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22187_ _03834_ _03836_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__nor2_1
XFILLER_0_218_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_217_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21138_ _02866_ _02881_ _02888_ _02880_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13960_ _06664_ _06679_ VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__nand2_1
X_21069_ _02745_ _02786_ _02744_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__o21ba_1
X_12911_ _05713_ _05714_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_1405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13891_ _06626_ _06620_ VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15630_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[4\] _08219_ _08220_
+ VGND VGND VPWR VPWR _08248_ sky130_fd_sc_hd__a21boi_2
X_12842_ _05647_ _05648_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__nor2_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15561_ net1027 _06660_ _08182_ _08166_ VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__o211a_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _05507_ _05581_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__or2_1
XFILLER_0_185_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _09842_ _09843_ VGND VGND VPWR VPWR _09844_ sky130_fd_sc_hd__nor2_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _07087_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[5\] _07060_
+ _07065_ VGND VGND VPWR VPWR _07205_ sky130_fd_sc_hd__and4_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18280_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[6\] _10747_ _08307_
+ VGND VGND VPWR VPWR _10748_ sky130_fd_sc_hd__mux2_1
X_15492_ _08116_ _08131_ VGND VGND VPWR VPWR _08132_ sky130_fd_sc_hd__nor2_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17231_ _09733_ _09734_ VGND VGND VPWR VPWR _09778_ sky130_fd_sc_hd__nand2_1
X_14443_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[4\] _07136_ _07137_
+ VGND VGND VPWR VPWR _07138_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17162_ _09699_ _09686_ _09711_ VGND VGND VPWR VPWR _09712_ sky130_fd_sc_hd__a21oi_1
X_14374_ top_inst.skew_buff_inst.row\[1\].output_reg\[4\] top_inst.axis_in_inst.inbuf_bus\[12\]
+ net207 VGND VGND VPWR VPWR _07077_ sky130_fd_sc_hd__mux2_4
XFILLER_0_80_942 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16113_ net1068 _08183_ _08702_ _08692_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13325_ _06099_ VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17093_ _09642_ _09643_ _09644_ VGND VGND VPWR VPWR _09645_ sky130_fd_sc_hd__nand3_1
XFILLER_0_150_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16044_ _08633_ _08650_ VGND VGND VPWR VPWR _08651_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13256_ _05992_ _05994_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_1287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12207_ top_inst.axis_out_inst.out_buff_data\[29\] _05129_ VGND VGND VPWR VPWR _05133_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_62_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13187_ _05886_ _05965_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__and2_1
XFILLER_0_202_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19803_ _01614_ _01615_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__or2b_1
X_12138_ net854 _05084_ _05093_ _05088_ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17995_ _10040_ _10300_ _10419_ _10459_ VGND VGND VPWR VPWR _10498_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_1186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16946_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[9\] _09459_ _09417_
+ VGND VGND VPWR VPWR _09501_ sky130_fd_sc_hd__a21o_1
X_19734_ _01561_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__clkbuf_4
X_12069_ net447 _05045_ _05054_ _05049_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_1_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_193_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19665_ _01492_ _01493_ _01494_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__and3_1
XFILLER_0_223_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16877_ _09431_ _09432_ _09433_ VGND VGND VPWR VPWR _09434_ sky130_fd_sc_hd__nand3_1
XFILLER_0_189_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18616_ _11065_ _11068_ VGND VGND VPWR VPWR _11075_ sky130_fd_sc_hd__or2_1
XFILLER_0_204_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15828_ _08439_ _08440_ VGND VGND VPWR VPWR _08441_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_205_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19596_ _01426_ _01427_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_231_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18547_ _10969_ _11007_ VGND VGND VPWR VPWR _11008_ sky130_fd_sc_hd__nor2_1
XFILLER_0_220_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15759_ _08371_ _08373_ VGND VGND VPWR VPWR _08374_ sky130_fd_sc_hd__nor2_4
XFILLER_0_73_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18478_ _10939_ _10940_ VGND VGND VPWR VPWR _10941_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_213_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17429_ _09965_ _09966_ VGND VGND VPWR VPWR _09967_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20440_ _02185_ _02202_ _02203_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__nor3_1
XFILLER_0_172_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_209_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20371_ _02155_ _02156_ _02148_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__a21o_1
XFILLER_0_141_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22110_ _03777_ _03801_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23090_ net25 _04600_ _04642_ _04643_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22041_ net1103 _09804_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__or2_1
XTAP_6409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_239_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_1163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23992_ clknet_leaf_79_clk _00525_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_199_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22943_ net732 _04548_ _04559_ _04551_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22874_ net296 _04517_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24613_ clknet_leaf_21_clk _01146_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_190_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21825_ _03486_ _03506_ _03545_ _03542_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__and4_1
XFILLER_0_167_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24544_ clknet_leaf_100_clk _01077_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dfxtp_2
X_21756_ _03456_ _03471_ _03480_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_231_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20707_ _02457_ _02485_ VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24475_ clknet_leaf_37_clk _01008_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_21687_ _03412_ _03413_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23426_ top_inst.axis_out_inst.out_buff_data\[102\] _04596_ VGND VGND VPWR VPWR _04834_
+ sky130_fd_sc_hd__or2_1
X_20638_ _02390_ _02418_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__xor2_2
XFILLER_0_164_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23357_ net42 _04792_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20569_ _02343_ _02345_ _02350_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13110_ top_inst.grid_inst.data_path_wires\[1\]\[0\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__or2b_1
X_22308_ _03986_ _03994_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__xnor2_2
X_14090_ _05632_ _06805_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23288_ net136 _04753_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13041_ _05734_ _05768_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__nand2_1
X_22239_ net817 _09804_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16800_ _08831_ _09358_ VGND VGND VPWR VPWR _09359_ sky130_fd_sc_hd__and2_1
XFILLER_0_218_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17780_ _10286_ _10287_ VGND VGND VPWR VPWR _10288_ sky130_fd_sc_hd__nor2_1
XFILLER_0_206_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_205_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14992_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[0\] _06660_ _07647_
+ _07643_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_1263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16731_ _05327_ VGND VGND VPWR VPWR _09292_ sky130_fd_sc_hd__buf_8
XFILLER_0_205_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13943_ _06656_ _06661_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19450_ net218 _01236_ _01283_ _01284_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_242_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16662_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[1\] _09224_ _09225_
+ VGND VGND VPWR VPWR _09226_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13874_ _06612_ _06613_ VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18401_ _10864_ _10865_ VGND VGND VPWR VPWR _10866_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15613_ _08207_ _08208_ _08231_ VGND VGND VPWR VPWR _08232_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_213_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19381_ _01210_ _01211_ _01217_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__and3_1
X_12825_ _04867_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_243_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16593_ _09143_ _09144_ _09141_ VGND VGND VPWR VPWR _09168_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18332_ _10589_ _10606_ _10608_ _10604_ VGND VGND VPWR VPWR _10798_ sky130_fd_sc_hd__nand4_2
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15544_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _08169_ sky130_fd_sc_hd__buf_2
X_12756_ _05304_ _05528_ _05292_ _05302_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__a22o_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18263_ _10606_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[2\] _10728_
+ _10729_ VGND VGND VPWR VPWR _10731_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15475_ _08088_ _08090_ _08114_ _08115_ VGND VGND VPWR VPWR _08116_ sky130_fd_sc_hd__and4bb_1
X_12687_ _05293_ _05288_ _05292_ _05297_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__and4_1
X_17214_ _09749_ _09750_ _09760_ VGND VGND VPWR VPWR _09762_ sky130_fd_sc_hd__and3_1
XFILLER_0_170_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14426_ _07119_ _07120_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[3\]
+ VGND VGND VPWR VPWR _07122_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_167_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18194_ top_inst.grid_inst.data_path_wires\[12\]\[3\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[12\]\[4\]
+ VGND VGND VPWR VPWR _10664_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17145_ _09695_ VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14357_ _05290_ _07061_ _07063_ _06684_ VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold707 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[24\] VGND
+ VGND VPWR VPWR net889 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ _05751_ _05770_ _06082_ _05748_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_122_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold718 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[24\] VGND
+ VGND VPWR VPWR net900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17076_ _09459_ VGND VGND VPWR VPWR _09628_ sky130_fd_sc_hd__clkbuf_4
Xhold729 top_inst.deskew_buff_inst.col_input\[6\] VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14288_ _06963_ top_inst.grid_inst.data_path_wires\[3\]\[6\] _06997_ VGND VGND VPWR
+ VPWR _06998_ sky130_fd_sc_hd__o21a_1
X_16027_ _08633_ _08634_ VGND VGND VPWR VPWR _08635_ sky130_fd_sc_hd__and2_1
X_13239_ top_inst.grid_inst.data_path_wires\[1\]\[7\] _05765_ _05763_ VGND VGND VPWR
+ VPWR _06016_ sky130_fd_sc_hd__and3_2
XFILLER_0_126_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_204_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1016 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17978_ _10450_ _10481_ VGND VGND VPWR VPWR _10482_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16929_ _09439_ _09458_ _09483_ _09484_ VGND VGND VPWR VPWR _09485_ sky130_fd_sc_hd__a211o_1
X_19717_ _01531_ _01544_ _01545_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__and3_1
XFILLER_0_237_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19648_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[10\] _01395_ _01396_
+ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19579_ _01408_ _01409_ _01407_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21610_ _03269_ _03276_ _03307_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_215_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22590_ _04137_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21541_ net839 _02638_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24260_ clknet_leaf_110_clk _00793_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21472_ _03201_ _03204_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_1307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23211_ _04686_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__buf_2
XFILLER_0_44_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20423_ _02206_ _02207_ _02139_ _02142_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__a211o_1
X_24191_ clknet_leaf_47_clk _00724_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23142_ net60 _04672_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__or2_1
X_20354_ _02139_ _02140_ _02102_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__o21a_1
XFILLER_0_222_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23073_ net16 _04628_ _04634_ _04632_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20285_ _02074_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__clkbuf_1
XTAP_6206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22024_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[1\] _03718_ _03719_
+ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__nand3_1
XTAP_6239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold78 top_inst.deskew_buff_inst.col_input\[117\] VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23975_ clknet_leaf_87_clk _00508_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_192_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold89 _00119_ VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_242_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22926_ _04868_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_196_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22857_ _02706_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12610_ _05378_ _05381_ _05379_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__a21bo_1
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21808_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[23\] _03376_ VGND
+ VGND VPWR VPWR _03530_ sky130_fd_sc_hd__xnor2_1
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13590_ _06336_ _06337_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22788_ _04438_ _04456_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12541_ _05342_ _05355_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__nor2_1
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24527_ clknet_leaf_128_clk _01060_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21739_ _03436_ _03445_ _03463_ _01984_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__a31o_1
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15260_ _06848_ _07905_ _07906_ _07643_ VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12472_ _05293_ _05294_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__or2_1
X_24458_ clknet_leaf_52_clk _00991_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14211_ _06364_ _06923_ VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__and2_1
X_23409_ net68 _04658_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15191_ _07746_ _07785_ _07838_ VGND VGND VPWR VPWR _07839_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_85_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24389_ clknet_leaf_38_clk _00922_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[0\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_14142_ _06854_ _06855_ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14073_ _06787_ _06788_ VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__or2_1
X_18950_ _11370_ _11372_ VGND VGND VPWR VPWR _11373_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13024_ _05804_ _05805_ _05790_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__a21oi_1
X_17901_ _10393_ _10366_ VGND VGND VPWR VPWR _10406_ sky130_fd_sc_hd__or2b_1
XFILLER_0_219_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18881_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[7\] _11304_ VGND
+ VGND VPWR VPWR _11305_ sky130_fd_sc_hd__xor2_2
XTAP_6740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17832_ _10035_ _10054_ VGND VGND VPWR VPWR _10339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17763_ _10184_ _10223_ VGND VGND VPWR VPWR _10272_ sky130_fd_sc_hd__nor2_1
XFILLER_0_206_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14975_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _07635_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16714_ _09193_ _09188_ _09202_ _09206_ VGND VGND VPWR VPWR _09275_ sky130_fd_sc_hd__nand4_1
X_19502_ net241 _01331_ _01332_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__or3_4
XFILLER_0_215_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13926_ _06630_ _06647_ _06651_ _06639_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17694_ _10170_ _10175_ VGND VGND VPWR VPWR _10204_ sky130_fd_sc_hd__and2_1
XFILLER_0_159_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19433_ _01261_ net232 _01267_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__nand3_2
XFILLER_0_202_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16645_ _09185_ _09210_ _09212_ _09184_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_1076 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13857_ _06596_ _06587_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__and2b_1
XFILLER_0_230_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_664 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12808_ _05507_ _05615_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19364_ _01201_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16576_ _09007_ _09121_ VGND VGND VPWR VPWR _09151_ sky130_fd_sc_hd__and2b_1
XFILLER_0_130_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13788_ _06528_ _06530_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18315_ _10744_ _10746_ _10743_ VGND VGND VPWR VPWR _10782_ sky130_fd_sc_hd__o21bai_2
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15527_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _08157_ sky130_fd_sc_hd__clkbuf_4
X_12739_ _05547_ _05548_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__and2_1
X_19295_ top_inst.skew_buff_inst.row\[3\].output_reg\[4\] top_inst.axis_in_inst.inbuf_bus\[28\]
+ net34 VGND VGND VPWR VPWR _11695_ sky130_fd_sc_hd__mux2_4
XFILLER_0_155_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18246_ _10691_ _10697_ VGND VGND VPWR VPWR _10714_ sky130_fd_sc_hd__or2b_1
XFILLER_0_199_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15458_ _08099_ VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14409_ _07103_ _07104_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[2\]
+ VGND VGND VPWR VPWR _07106_ sky130_fd_sc_hd__a21o_1
XFILLER_0_163_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18177_ _10581_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[0\]
+ _10585_ VGND VGND VPWR VPWR _10648_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15389_ _07622_ _07824_ _08031_ VGND VGND VPWR VPWR _08032_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17128_ _09673_ _09676_ _09677_ _09678_ VGND VGND VPWR VPWR _09679_ sky130_fd_sc_hd__a211o_1
Xhold504 top_inst.axis_out_inst.out_buff_data\[5\] VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold515 top_inst.axis_out_inst.out_buff_data\[105\] VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold526 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[7\] VGND VGND
+ VPWR VPWR net708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold537 _00962_ VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold548 top_inst.axis_out_inst.out_buff_data\[62\] VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__dlygate4sd3_1
X_17059_ _09562_ _09563_ _09564_ _09567_ VGND VGND VPWR VPWR _09612_ sky130_fd_sc_hd__a31o_1
XFILLER_0_180_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold559 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[5\] VGND
+ VGND VPWR VPWR net741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20070_ _01864_ _01867_ _01884_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__o21ai_2
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20972_ _02727_ _02728_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__nand2_1
X_23760_ clknet_leaf_123_clk net336 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22711_ net441 _09804_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23691_ clknet_leaf_120_clk _00224_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22642_ _04287_ _04294_ _04313_ _04267_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22573_ _04231_ _04250_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24312_ clknet_leaf_1_clk _00845_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[87\]
+ sky130_fd_sc_hd__dfxtp_1
X_21524_ _03253_ _03256_ VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21455_ _03154_ _03189_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__xor2_2
X_24243_ clknet_leaf_116_clk _00776_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20406_ top_inst.grid_inst.data_path_wires\[16\]\[4\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[3\]
+ _02051_ top_inst.grid_inst.data_path_wires\[16\]\[5\] VGND VGND VPWR VPWR _02192_
+ sky130_fd_sc_hd__a22o_1
X_24174_ clknet_leaf_23_clk _00707_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21386_ _03080_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_189_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23125_ net463 _04656_ _04664_ _04662_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__o211a_1
X_20337_ _02100_ _02101_ _02124_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__a21o_1
XTAP_6003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput46 net46 VGND VGND VPWR VPWR output_tdata[107] sky130_fd_sc_hd__buf_2
XFILLER_0_101_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23056_ net8 _04615_ _04624_ _04619_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__o211a_1
Xoutput57 net57 VGND VGND VPWR VPWR output_tdata[117] sky130_fd_sc_hd__clkbuf_4
XTAP_6025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput68 net68 VGND VGND VPWR VPWR output_tdata[127] sky130_fd_sc_hd__buf_2
X_20268_ _02057_ _02055_ _02038_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_101_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput79 net79 VGND VGND VPWR VPWR output_tdata[21] sky130_fd_sc_hd__clkbuf_4
XTAP_6047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22007_ _03707_ _05275_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__or2_1
XTAP_6069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20199_ _04858_ _11705_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__or2_2
XTAP_5346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14760_ _07407_ _07406_ VGND VGND VPWR VPWR _07447_ sky130_fd_sc_hd__or2b_1
XTAP_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ top_inst.axis_out_inst.out_buff_data\[56\] _04996_ VGND VGND VPWR VPWR _04999_
+ sky130_fd_sc_hd__or2_1
X_23958_ clknet_leaf_89_clk _00491_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13711_ _06411_ _06414_ _06412_ VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_19_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22909_ top_inst.skew_buff_inst.row\[2\].output_reg\[2\] _04530_ VGND VGND VPWR VPWR
+ _04540_ sky130_fd_sc_hd__or2_1
XTAP_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14691_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[7\] _07333_ _07078_
+ _07087_ VGND VGND VPWR VPWR _07380_ sky130_fd_sc_hd__a22o_1
XTAP_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23889_ clknet_leaf_63_clk _00422_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16430_ _08876_ top_inst.grid_inst.data_path_wires\[8\]\[4\] top_inst.grid_inst.data_path_wires\[8\]\[5\]
+ _08697_ VGND VGND VPWR VPWR _09009_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_39_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13642_ _06384_ _06345_ _06387_ _06388_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__o211a_1
XFILLER_0_224_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16361_ _08940_ _08941_ VGND VGND VPWR VPWR _08942_ sky130_fd_sc_hd__nor2_1
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13573_ _06289_ _06285_ _06320_ _06321_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__a211oi_2
X_18100_ _10029_ _10584_ _10586_ _10448_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15312_ top_inst.grid_inst.data_path_wires\[6\]\[4\] VGND VGND VPWR VPWR _07957_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_81_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12524_ _05338_ _05339_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__nor2_1
X_19080_ _11498_ _11499_ VGND VGND VPWR VPWR _11500_ sky130_fd_sc_hd__and2_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[7\] _08862_ VGND
+ VGND VPWR VPWR _08874_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18031_ _10531_ _10532_ VGND VGND VPWR VPWR _10533_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_164_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15243_ _07833_ _07835_ _07888_ VGND VGND VPWR VPWR _07890_ sky130_fd_sc_hd__and3_1
X_12455_ _05280_ _05276_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15174_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[7\] _07810_ VGND
+ VGND VPWR VPWR _07822_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12386_ _05142_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_105_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14125_ _06795_ _06797_ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__or2b_1
XFILLER_0_22_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19982_ _01779_ _01781_ _01799_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__a21o_1
XFILLER_0_162_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_674 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14056_ _06770_ _06771_ VGND VGND VPWR VPWR _06772_ sky130_fd_sc_hd__xnor2_2
X_18933_ _11161_ _11135_ _11317_ _11355_ VGND VGND VPWR VPWR _11356_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_219_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13007_ _05789_ _05790_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18864_ _11286_ _11287_ _11258_ _11259_ VGND VGND VPWR VPWR _11289_ sky130_fd_sc_hd__o211ai_1
XTAP_6570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17815_ net1016 _09266_ _10321_ _10322_ _09886_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__o221a_1
X_18795_ _11216_ _11221_ VGND VGND VPWR VPWR _11222_ sky130_fd_sc_hd__xnor2_2
XTAP_5880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17746_ _10169_ _10214_ VGND VGND VPWR VPWR _10255_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14958_ _07622_ _07611_ _07623_ _07618_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13909_ _06618_ _06204_ _06638_ _06639_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17677_ _10186_ _10187_ VGND VGND VPWR VPWR _10188_ sky130_fd_sc_hd__nor2_1
X_14889_ _07558_ _07572_ VGND VGND VPWR VPWR _07573_ sky130_fd_sc_hd__xor2_2
XFILLER_0_203_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_230_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16628_ _05772_ VGND VGND VPWR VPWR _09199_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19416_ _01218_ _01219_ _01220_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_187_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16559_ _09133_ _09134_ VGND VGND VPWR VPWR _09135_ sky130_fd_sc_hd__nand2_1
X_19347_ _11693_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[2\] net243
+ _11682_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__nand4_1
XFILLER_0_31_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1069 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19278_ top_inst.skew_buff_inst.row\[3\].output_reg\[1\] top_inst.axis_in_inst.inbuf_bus\[25\]
+ net188 VGND VGND VPWR VPWR _11681_ sky130_fd_sc_hd__mux2_4
XFILLER_0_116_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18229_ _10691_ _10697_ VGND VGND VPWR VPWR _10698_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21240_ _02971_ _02979_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__xor2_2
XFILLER_0_241_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold301 top_inst.deskew_buff_inst.col_input\[14\] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold312 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[3\] VGND
+ VGND VPWR VPWR net494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[15\] VGND
+ VGND VPWR VPWR net505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _00277_ VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21171_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[2\] _02913_ VGND
+ VGND VPWR VPWR _02914_ sky130_fd_sc_hd__xor2_1
Xhold345 _00192_ VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[14\] VGND
+ VGND VPWR VPWR net538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[13\] VGND
+ VGND VPWR VPWR net549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20122_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[28\] _01761_ _01762_
+ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__a21o_1
XFILLER_0_141_1143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold378 _00133_ VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 _00021_ VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20053_ _01783_ _01850_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23812_ clknet_leaf_72_clk _00345_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23743_ clknet_leaf_122_clk _00276_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20955_ _02643_ _02723_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__xnor2_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23674_ clknet_leaf_116_clk net847 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20886_ _02656_ _02657_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_1302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22625_ _04284_ _04301_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22556_ _04208_ _04211_ _04234_ _06734_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21507_ _03225_ _03223_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__or2b_1
XFILLER_0_161_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22487_ _04164_ _04168_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12240_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[11\] _05143_
+ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__or2_1
X_24226_ clknet_leaf_112_clk _00759_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[16\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21438_ top_inst.grid_inst.data_path_wires\[17\]\[3\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12171_ net359 _05102_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__or2_1
X_24157_ clknet_leaf_17_clk _00690_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_20_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21369_ _03058_ _03035_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__or2b_1
XFILLER_0_124_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23108_ net331 _10541_ _04652_ _04643_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24088_ clknet_leaf_87_clk _00621_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold890 top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[3\] VGND VGND
+ VPWR VPWR net1072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15930_ _08500_ _08499_ VGND VGND VPWR VPWR _08541_ sky130_fd_sc_hd__or2b_1
X_23039_ net32 _04601_ _04614_ _04606_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__o211a_1
XTAP_5110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15861_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[10\] _08066_ _08472_
+ _08473_ VGND VGND VPWR VPWR _08474_ sky130_fd_sc_hd__a22o_1
XTAP_5165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _10111_ _10112_ VGND VGND VPWR VPWR _10113_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_235_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14812_ _07241_ _07086_ _07496_ VGND VGND VPWR VPWR _07498_ sky130_fd_sc_hd__o21ai_1
XTAP_5198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18580_ _10960_ _10998_ _11036_ _11039_ _11035_ VGND VGND VPWR VPWR _11040_ sky130_fd_sc_hd__a32o_1
XFILLER_0_203_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15792_ top_inst.grid_inst.data_path_wires\[7\]\[6\] top_inst.grid_inst.data_path_wires\[7\]\[5\]
+ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _08406_ sky130_fd_sc_hd__and4_1
XFILLER_0_99_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_235_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _10052_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14743_ _07428_ _07429_ _07430_ VGND VGND VPWR VPWR _07431_ sky130_fd_sc_hd__nand3_1
XTAP_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ net876 _04977_ _04988_ _04981_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17462_ _09978_ _09993_ _09997_ VGND VGND VPWR VPWR _09998_ sky130_fd_sc_hd__o21a_1
X_14674_ _07319_ _07323_ _07322_ VGND VGND VPWR VPWR _07363_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_196_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11886_ net878 _04938_ _04949_ _04942_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16413_ _08920_ _08914_ _08954_ VGND VGND VPWR VPWR _08993_ sky130_fd_sc_hd__a21oi_1
X_19201_ _11177_ _11616_ _11617_ _11160_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13625_ _06330_ _06331_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17393_ _09892_ _09930_ _09931_ VGND VGND VPWR VPWR _09932_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19132_ _11512_ _11518_ _11516_ VGND VGND VPWR VPWR _11550_ sky130_fd_sc_hd__a21o_1
XFILLER_0_171_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16344_ _08923_ _08924_ VGND VGND VPWR VPWR _08925_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13556_ _06265_ _06268_ _06266_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_15_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19063_ _11481_ VGND VGND VPWR VPWR _11483_ sky130_fd_sc_hd__inv_2
X_12507_ _05324_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__clkbuf_16
X_16275_ _08807_ _08813_ VGND VGND VPWR VPWR _08858_ sky130_fd_sc_hd__or2b_1
X_13487_ _06227_ _06237_ _06238_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__nor3_1
X_18014_ _10486_ _10516_ VGND VGND VPWR VPWR _10517_ sky130_fd_sc_hd__xor2_1
X_15226_ _07615_ _07637_ VGND VGND VPWR VPWR _07873_ sky130_fd_sc_hd__nand2_1
X_12438_ net34 VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__buf_8
XFILLER_0_113_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15157_ _07755_ _07762_ VGND VGND VPWR VPWR _07806_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12369_ net848 _05217_ _05225_ _05221_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_238_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14108_ _06820_ _06822_ VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19965_ _01783_ _01769_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__nor2_1
X_15088_ _07117_ _07738_ VGND VGND VPWR VPWR _07739_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14039_ _06749_ _06755_ VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__xnor2_2
X_18916_ top_inst.grid_inst.data_path_wires\[13\]\[7\] _11152_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _11339_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19896_ _01704_ _01707_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__or2b_1
XFILLER_0_219_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18847_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[5\] _11132_ top_inst.grid_inst.data_path_wires\[13\]\[0\]
+ _11164_ VGND VGND VPWR VPWR _11272_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_59_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18778_ _11203_ _11204_ _11190_ VGND VGND VPWR VPWR _11206_ sky130_fd_sc_hd__a21o_1
XFILLER_0_222_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17729_ _10233_ _10237_ VGND VGND VPWR VPWR _10238_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20740_ _02364_ _02440_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__nand2_2
XFILLER_0_148_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20671_ _02416_ _02450_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22410_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[12\] _03937_ _03938_
+ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23390_ net58 _04805_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__or2_1
XFILLER_0_169_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22341_ top_inst.grid_inst.data_path_wires\[18\]\[4\] _03713_ VGND VGND VPWR VPWR
+ _04027_ sky130_fd_sc_hd__and2b_1
XFILLER_0_171_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22272_ _03951_ _03959_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24011_ clknet_leaf_47_clk _00544_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21223_ _02939_ _02958_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__nor2_1
Xhold120 top_inst.deskew_buff_inst.col_input\[102\] VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold131 top_inst.deskew_buff_inst.col_input\[67\] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold142 _00182_ VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[30\] VGND
+ VGND VPWR VPWR net335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[16\] VGND
+ VGND VPWR VPWR net346 sky130_fd_sc_hd__dlygate4sd3_1
X_21154_ _02862_ _02883_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__and3_1
Xhold175 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[10\] VGND
+ VGND VPWR VPWR net357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold186 _00016_ VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 top_inst.axis_out_inst.out_buff_data\[24\] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20105_ _01563_ _01917_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21085_ _02821_ _02825_ _02836_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__o21a_1
XFILLER_0_186_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20036_ _01850_ _01851_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__xor2_1
XFILLER_0_232_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21987_ _03693_ _03691_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _04861_ _04856_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__nor2_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23726_ clknet_leaf_121_clk _00259_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ _01819_ _02704_ _02705_ _02707_ VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__o211a_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23657_ clknet_leaf_132_clk net366 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_20869_ _02632_ _02636_ _02640_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_187_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13410_ top_inst.grid_inst.data_path_wires\[2\]\[0\] VGND VGND VPWR VPWR _06181_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22608_ _04268_ _04267_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14390_ _07089_ VGND VGND VPWR VPWR _07090_ sky130_fd_sc_hd__buf_4
XFILLER_0_193_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23588_ clknet_leaf_106_clk net269 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13341_ top_inst.grid_inst.data_path_wires\[1\]\[7\] _05770_ VGND VGND VPWR VPWR
+ _06115_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22539_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[17\] _04163_ VGND
+ VGND VPWR VPWR _04219_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16060_ _08664_ _08140_ VGND VGND VPWR VPWR _08665_ sky130_fd_sc_hd__or2_1
X_13272_ _06046_ _06047_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15011_ _07653_ _07664_ VGND VGND VPWR VPWR _07665_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12223_ _04863_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__clkbuf_4
X_24209_ clknet_leaf_118_clk _00742_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_972 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12154_ top_inst.axis_out_inst.out_buff_data\[6\] _05102_ VGND VGND VPWR VPWR _05103_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_102_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_1346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_236_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19750_ _01575_ _01576_ _01488_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_235_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16962_ _09513_ _09514_ _09515_ VGND VGND VPWR VPWR _09517_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_1212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12085_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[8\] _05063_
+ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__or2_1
X_18701_ top_inst.grid_inst.data_path_wires\[13\]\[5\] VGND VGND VPWR VPWR _11143_
+ sky130_fd_sc_hd__clkbuf_4
X_15913_ _08522_ _08523_ VGND VGND VPWR VPWR _08524_ sky130_fd_sc_hd__xor2_1
XFILLER_0_99_1380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16893_ _09409_ _09449_ VGND VGND VPWR VPWR _09450_ sky130_fd_sc_hd__xor2_1
X_19681_ net1116 _01510_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_194_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15844_ _08453_ _08456_ VGND VGND VPWR VPWR _08457_ sky130_fd_sc_hd__xor2_1
X_18632_ _11088_ _11089_ VGND VGND VPWR VPWR _11091_ sky130_fd_sc_hd__nand2_1
XTAP_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15775_ _08387_ _08389_ VGND VGND VPWR VPWR _08390_ sky130_fd_sc_hd__xnor2_1
X_18563_ _11012_ _10984_ _11023_ VGND VGND VPWR VPWR _11024_ sky130_fd_sc_hd__a21o_1
XFILLER_0_235_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12987_ _05753_ _05756_ _05774_ _05767_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__o211a_1
XTAP_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _07412_ _07413_ VGND VGND VPWR VPWR _07414_ sky130_fd_sc_hd__nor2_2
X_17514_ top_inst.grid_inst.data_path_wires\[11\]\[7\] VGND VGND VPWR VPWR _10040_
+ sky130_fd_sc_hd__buf_4
XTAP_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18494_ _05633_ VGND VGND VPWR VPWR _10957_ sky130_fd_sc_hd__buf_4
XFILLER_0_115_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11938_ net613 _04969_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__or2_1
XFILLER_0_197_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17445_ _09952_ _09962_ _09981_ VGND VGND VPWR VPWR _09982_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_185_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14657_ _07284_ _07301_ VGND VGND VPWR VPWR _07347_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11869_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[12\] _04930_
+ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13608_ _06313_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__inv_2
X_17376_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[24\] _09628_ _09629_
+ VGND VGND VPWR VPWR _09916_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14588_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[0\]
+ _07089_ VGND VGND VPWR VPWR _07279_ sky130_fd_sc_hd__and3_1
XFILLER_0_166_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16327_ _08846_ _08853_ _08851_ VGND VGND VPWR VPWR _08909_ sky130_fd_sc_hd__a21oi_1
X_19115_ _11531_ _11533_ VGND VGND VPWR VPWR _11534_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13539_ _06288_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19046_ _11177_ _11465_ _11466_ _11160_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16258_ _08673_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[2\] _08839_
+ _08840_ VGND VGND VPWR VPWR _08841_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15209_ _07794_ _07801_ _07799_ VGND VGND VPWR VPWR _07857_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_23_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16189_ _08673_ top_inst.grid_inst.data_path_wires\[8\]\[4\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[1\]
+ _08682_ VGND VGND VPWR VPWR _08774_ sky130_fd_sc_hd__nand4_1
XFILLER_0_3_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19948_ _01766_ _01767_ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__nor2_1
XFILLER_0_177_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19879_ _01611_ _01688_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__or2_2
XFILLER_0_156_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21910_ net682 _03528_ _03626_ _03627_ _02962_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__o221a_1
X_22890_ net655 _04517_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21841_ _03554_ _03561_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_214_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24560_ clknet_leaf_134_clk _01093_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_77_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21772_ _03491_ _03495_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_172_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23511_ clknet_leaf_137_clk _00044_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_20723_ _02469_ _02500_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__xnor2_1
X_24491_ clknet_leaf_109_clk _01024_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_188_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23442_ top_inst.axis_out_inst.out_buff_data\[109\] _04835_ VGND VGND VPWR VPWR _04843_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_18_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20654_ _02432_ _02433_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_190_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23373_ net50 _04805_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__or2_1
X_20585_ _01999_ _02020_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22324_ _03311_ _04010_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22255_ _03941_ _03942_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1008 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21206_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[4\] _02946_ VGND
+ VGND VPWR VPWR _02947_ sky130_fd_sc_hd__xor2_2
X_22186_ _03848_ _03875_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_1311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21137_ _02887_ _02021_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__or2_1
XFILLER_0_217_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21068_ _02830_ _02831_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__nand2_1
XFILLER_0_217_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12910_ _05713_ _05714_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__or2_1
X_20019_ _01834_ _01835_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__and2_1
XFILLER_0_232_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13890_ top_inst.grid_inst.data_path_wires\[3\]\[3\] VGND VGND VPWR VPWR _06626_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12841_ _05645_ _05646_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__and2_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _08179_ _08180_ _08181_ VGND VGND VPWR VPWR _08182_ sky130_fd_sc_hd__o21ai_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12772_ _05535_ _05538_ _05536_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__o21ba_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _07087_ _07060_ _07065_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[5\]
+ VGND VGND VPWR VPWR _07204_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_185_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23709_ clknet_leaf_124_clk _00242_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15491_ _08125_ _08130_ VGND VGND VPWR VPWR _08131_ sky130_fd_sc_hd__xnor2_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _09770_ _09776_ VGND VGND VPWR VPWR _09777_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_182_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14442_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[0\]
+ _07072_ _07077_ VGND VGND VPWR VPWR _07137_ sky130_fd_sc_hd__nand4_1
XFILLER_0_166_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17161_ _09701_ _09710_ VGND VGND VPWR VPWR _09711_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14373_ _05290_ _07073_ _07076_ _06684_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16112_ _08700_ _08701_ _08181_ VGND VGND VPWR VPWR _08702_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13324_ _06097_ _06098_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__nand2_2
XFILLER_0_243_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17092_ _09553_ _09603_ _09602_ VGND VGND VPWR VPWR _09644_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_162_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16043_ _08636_ _08637_ _08649_ VGND VGND VPWR VPWR _08650_ sky130_fd_sc_hd__o21a_1
X_13255_ _05989_ _06031_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_161_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12206_ net308 _05123_ _05132_ _05128_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__o211a_1
X_13186_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[8\] _05354_ _05963_
+ _05964_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__a22o_1
XFILLER_0_209_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19802_ _01597_ _01619_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12137_ net722 _05089_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__or2_1
XFILLER_0_236_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17994_ _10495_ _10496_ VGND VGND VPWR VPWR _10497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19733_ _01528_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__clkbuf_4
X_16945_ _09464_ _09481_ _09482_ VGND VGND VPWR VPWR _09500_ sky130_fd_sc_hd__nand3_2
X_12068_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[1\] _05050_
+ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__or2_1
XFILLER_0_236_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19664_ _01445_ _01447_ _01446_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__a21bo_1
X_16876_ _09376_ _09379_ _09378_ VGND VGND VPWR VPWR _09433_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_172_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18615_ _11040_ _11070_ _11073_ VGND VGND VPWR VPWR _11074_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_220_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ _08147_ _08167_ VGND VGND VPWR VPWR _08440_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19595_ _01349_ _01380_ _01378_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__a21o_1
XTAP_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18546_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[13\] _10923_ VGND
+ VGND VPWR VPWR _11007_ sky130_fd_sc_hd__xnor2_1
X_15758_ _08372_ VGND VGND VPWR VPWR _08373_ sky130_fd_sc_hd__clkbuf_4
XTAP_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14709_ _07360_ _07396_ _07397_ VGND VGND VPWR VPWR _07398_ sky130_fd_sc_hd__or3_4
XFILLER_0_47_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18477_ _10896_ _10898_ _10897_ VGND VGND VPWR VPWR _10940_ sky130_fd_sc_hd__o21ba_1
X_15689_ _08304_ _08305_ VGND VGND VPWR VPWR _08306_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_200_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17428_ _09963_ _09964_ VGND VGND VPWR VPWR _09966_ sky130_fd_sc_hd__and2_1
XFILLER_0_172_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17359_ _09726_ _09877_ VGND VGND VPWR VPWR _09900_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20370_ _02148_ _02155_ _02156_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__nand3_1
XFILLER_0_28_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19029_ _11436_ _11437_ _11449_ VGND VGND VPWR VPWR _11450_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22040_ _03723_ _03734_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1085 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23991_ clknet_leaf_79_clk _00524_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22942_ net396 _04557_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__or2_1
XFILLER_0_214_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22873_ net387 _04509_ _04519_ _04511_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24612_ clknet_leaf_31_clk _01145_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_39_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21824_ _03524_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__inv_2
XFILLER_0_211_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24543_ clknet_leaf_130_clk _01076_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dfxtp_4
X_21755_ _03472_ _03479_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_210_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20706_ _02483_ _02484_ VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__xnor2_1
X_24474_ clknet_leaf_37_clk _01007_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21686_ _03412_ _03413_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23425_ net424 _04827_ _04833_ _04831_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20637_ _02416_ _02417_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23356_ net679 _04791_ _04796_ _04795_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20568_ _02311_ _02342_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22307_ _03991_ _03993_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__xor2_2
X_23287_ net757 _04752_ _04757_ _04756_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__o211a_1
X_20499_ top_inst.grid_inst.data_path_wires\[16\]\[3\] _02020_ VGND VGND VPWR VPWR
+ _02283_ sky130_fd_sc_hd__nand2_1
X_13040_ _05809_ _05814_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22238_ _03887_ _03926_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__xor2_1
XFILLER_0_218_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22169_ _03857_ _03858_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14991_ _07645_ _07646_ _05336_ VGND VGND VPWR VPWR _07647_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16730_ _09289_ _09290_ VGND VGND VPWR VPWR _09291_ sky130_fd_sc_hd__nor2_1
X_13942_ _06640_ _06622_ _06637_ _06624_ VGND VGND VPWR VPWR _06663_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16661_ _09194_ _09189_ _09187_ _09192_ VGND VGND VPWR VPWR _09225_ sky130_fd_sc_hd__nand4_1
XFILLER_0_57_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13873_ _06542_ _06595_ _06593_ VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_242_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18400_ _10847_ _10848_ _10863_ VGND VGND VPWR VPWR _10865_ sky130_fd_sc_hd__and3_1
X_15612_ _08202_ _08209_ VGND VGND VPWR VPWR _08231_ sky130_fd_sc_hd__or2_1
X_12824_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[11\] _05314_ _05631_
+ _05308_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16592_ _09137_ _09139_ _09166_ VGND VGND VPWR VPWR _09167_ sky130_fd_sc_hd__o21ba_1
X_19380_ _01215_ _01216_ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__and2_1
XFILLER_0_232_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15543_ _08147_ _07639_ _08168_ _08166_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__o211a_1
X_18331_ _10606_ _10608_ _10604_ _10589_ VGND VGND VPWR VPWR _10797_ sky130_fd_sc_hd__a22o_1
X_12755_ _05532_ _05533_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__or2_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18262_ _10728_ _10729_ _10606_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[2\]
+ VGND VGND VPWR VPWR _10730_ sky130_fd_sc_hd__and4bb_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _08112_ _08113_ VGND VGND VPWR VPWR _08115_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12686_ _05293_ _05292_ _05297_ _05288_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_182_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17213_ _09749_ _09750_ _09760_ VGND VGND VPWR VPWR _09761_ sky130_fd_sc_hd__a21oi_1
X_14425_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[3\] _07119_ _07120_
+ VGND VGND VPWR VPWR _07121_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18193_ _10663_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17144_ _09661_ _09694_ VGND VGND VPWR VPWR _09695_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14356_ _07062_ _06641_ VGND VGND VPWR VPWR _07063_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13307_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _06082_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold708 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[16\] VGND
+ VGND VPWR VPWR net890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17075_ _09590_ _09593_ _09626_ VGND VGND VPWR VPWR _09627_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold719 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[7\] VGND
+ VGND VPWR VPWR net901 sky130_fd_sc_hd__dlygate4sd3_1
X_14287_ top_inst.grid_inst.data_path_wires\[3\]\[7\] _06652_ VGND VGND VPWR VPWR
+ _06997_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_208_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16026_ _08628_ _08632_ VGND VGND VPWR VPWR _08634_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_243_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13238_ _06013_ _06014_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__xor2_1
XFILLER_0_228_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13169_ _05896_ _05898_ _05946_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__nand3_1
XFILLER_0_23_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17977_ _10479_ _10480_ VGND VGND VPWR VPWR _10481_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19716_ _01541_ _01542_ _01543_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__a21o_1
X_16928_ _09481_ _09482_ net200 VGND VGND VPWR VPWR _09484_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19647_ _01440_ _01456_ _01457_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__nand3_1
X_16859_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[0\]
+ _09217_ VGND VGND VPWR VPWR _09416_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19578_ _01407_ _01408_ _01409_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__nand3_1
XFILLER_0_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18529_ _10966_ _10990_ VGND VGND VPWR VPWR _10991_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21540_ _03238_ _03272_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21471_ _03201_ _03204_ VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23210_ _04684_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__clkbuf_4
X_20422_ _02139_ _02142_ _02206_ _02207_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_181_1319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24190_ clknet_leaf_48_clk _00723_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23141_ net440 _04671_ _04673_ _04662_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20353_ _02137_ _02138_ _02107_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23072_ net1110 _04629_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__or2_1
X_20284_ _11722_ _02073_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22023_ _03700_ _03682_ _03698_ _03680_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__nand4_2
XTAP_6229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23974_ clknet_leaf_87_clk _00507_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_242_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold79 _01174_ VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22925_ net643 _04543_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__or2_1
XFILLER_0_202_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_233_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22856_ net707 _04504_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21807_ _03494_ _03515_ _03513_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22787_ _04454_ _04455_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__xnor2_1
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12540_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[0\]
+ _05282_ _05287_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__and4_1
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24526_ clknet_leaf_128_clk _01059_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_213_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21738_ _03436_ _03445_ _03463_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24457_ clknet_leaf_58_clk _00990_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_12471_ _05275_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__buf_2
XFILLER_0_35_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21669_ _03336_ _03347_ _03365_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__a21bo_1
X_14210_ _06921_ _06922_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[10\]
+ _05327_ VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__a2bb2o_1
X_23408_ net623 _04655_ _04824_ _04819_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15190_ _07786_ _07789_ _07790_ VGND VGND VPWR VPWR _07838_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24388_ clknet_leaf_39_clk _00921_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14141_ _06807_ _06810_ _06808_ VGND VGND VPWR VPWR _06855_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23339_ net557 _04778_ _04786_ _04782_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_240_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14072_ _06784_ _06786_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13023_ _05790_ _05804_ _05805_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17900_ _10391_ _10392_ VGND VGND VPWR VPWR _10405_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18880_ _11302_ _11303_ VGND VGND VPWR VPWR _11304_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17831_ _10296_ _10337_ VGND VGND VPWR VPWR _10338_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_234_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_233_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17762_ _10269_ _10270_ VGND VGND VPWR VPWR _10271_ sky130_fd_sc_hd__nor2_1
X_14974_ _07613_ _06647_ _07634_ _07618_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__o211a_1
X_19501_ _01298_ _01333_ _01334_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__or3b_1
XFILLER_0_107_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16713_ _09193_ _09202_ _09206_ _09188_ VGND VGND VPWR VPWR _09274_ sky130_fd_sc_hd__a22o_1
X_13925_ _06650_ _06641_ VGND VGND VPWR VPWR _06651_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_1191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17693_ _10196_ _10202_ VGND VGND VPWR VPWR _10203_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19432_ _01264_ _01265_ _01239_ _01240_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_57_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16644_ _09211_ _09199_ VGND VGND VPWR VPWR _09212_ sky130_fd_sc_hd__or2_1
XFILLER_0_173_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13856_ _06587_ _06596_ VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12807_ _05538_ _05574_ _05575_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_202_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19363_ _11722_ _01200_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16575_ _09124_ _09131_ _09123_ VGND VGND VPWR VPWR _09150_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13787_ _06198_ _06212_ _06529_ VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18314_ _10741_ _10780_ VGND VGND VPWR VPWR _10781_ sky130_fd_sc_hd__xor2_1
X_12738_ _05507_ _05546_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15526_ _08135_ _07639_ _08156_ _08142_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19294_ _09185_ _11692_ _11694_ _11641_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15457_ _07117_ _08098_ VGND VGND VPWR VPWR _08099_ sky130_fd_sc_hd__and2_1
X_18245_ _10696_ _10692_ VGND VGND VPWR VPWR _10713_ sky130_fd_sc_hd__or2b_1
X_12669_ _05335_ _05478_ _05479_ _05480_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__a31o_1
XFILLER_0_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14408_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[2\] _07103_ _07104_
+ VGND VGND VPWR VPWR _07105_ sky130_fd_sc_hd__nand3_1
XFILLER_0_113_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15388_ _07624_ _07640_ VGND VGND VPWR VPWR _08031_ sky130_fd_sc_hd__nand2_1
X_18176_ _10644_ _10646_ VGND VGND VPWR VPWR _10647_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17127_ _09551_ _09552_ _09673_ VGND VGND VPWR VPWR _09678_ sky130_fd_sc_hd__a21oi_2
X_14339_ _05632_ _07047_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold505 top_inst.axis_out_inst.out_buff_data\[79\] VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[24\] VGND
+ VGND VPWR VPWR net698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 _00925_ VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold538 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[27\] VGND
+ VGND VPWR VPWR net720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17058_ _09609_ _09610_ VGND VGND VPWR VPWR _09611_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold549 top_inst.axis_out_inst.out_buff_data\[46\] VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16009_ _08585_ _08617_ VGND VGND VPWR VPWR _08618_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20971_ _01819_ _02738_ _02739_ _02707_ VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22710_ _04364_ _04382_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23690_ clknet_leaf_120_clk _00223_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22641_ _04315_ _04316_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22572_ _04231_ _04250_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24311_ clknet_leaf_2_clk _00844_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[86\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21523_ _03254_ _03255_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24242_ clknet_leaf_108_clk _00775_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_21454_ _03161_ _03188_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20405_ _02189_ _02190_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__xor2_2
XFILLER_0_107_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24173_ clknet_leaf_23_clk _00706_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_1235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21385_ _03076_ _03081_ _03120_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23124_ net99 _04659_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20336_ _02122_ _02123_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput47 net47 VGND VGND VPWR VPWR output_tdata[108] sky130_fd_sc_hd__clkbuf_4
Xoutput58 net58 VGND VGND VPWR VPWR output_tdata[118] sky130_fd_sc_hd__clkbuf_4
X_23055_ top_inst.axis_in_inst.inbuf_bus\[16\] _04616_ VGND VGND VPWR VPWR _04624_
+ sky130_fd_sc_hd__or2_1
XTAP_6015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput69 net69 VGND VGND VPWR VPWR output_tdata[12] sky130_fd_sc_hd__buf_2
XTAP_6026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20267_ _01993_ _02009_ _02052_ _02053_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__nand4_1
XTAP_6037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22006_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _03707_ sky130_fd_sc_hd__buf_2
XTAP_6059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20198_ top_inst.grid_inst.data_path_wires\[16\]\[6\] VGND VGND VPWR VPWR _02001_
+ sky130_fd_sc_hd__buf_4
XTAP_5336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_231_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23957_ clknet_leaf_91_clk _00490_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_4
X_11971_ net700 _04990_ _04998_ _04995_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__o211a_1
XTAP_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13710_ _06453_ _06454_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22908_ net769 _04535_ _04539_ _04537_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14690_ _07241_ _07242_ _07073_ _07378_ VGND VGND VPWR VPWR _07379_ sky130_fd_sc_hd__or4_1
XFILLER_0_169_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23888_ clknet_leaf_64_clk _00421_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13641_ _06335_ _06337_ _06386_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__nand3_1
XFILLER_0_211_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22839_ net406 _04496_ _04500_ _04498_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16360_ _08885_ _08887_ _08939_ VGND VGND VPWR VPWR _08941_ sky130_fd_sc_hd__and3_1
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13572_ _06315_ _06316_ _06319_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__o21a_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15311_ _07881_ _07955_ VGND VGND VPWR VPWR _07956_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_13_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12523_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[3\] top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[2\]
+ _05271_ _05278_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__and4_1
X_24509_ clknet_leaf_128_clk _01042_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dfxtp_4
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16291_ _08861_ _08860_ VGND VGND VPWR VPWR _08873_ sky130_fd_sc_hd__or2b_1
XFILLER_0_186_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15242_ _07833_ _07835_ _07888_ VGND VGND VPWR VPWR _07889_ sky130_fd_sc_hd__a21oi_1
X_18030_ _10495_ _10496_ _10506_ _10504_ VGND VGND VPWR VPWR _10532_ sky130_fd_sc_hd__a31o_1
XFILLER_0_240_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12454_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _05280_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_151_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15173_ _07809_ _07808_ VGND VGND VPWR VPWR _07821_ sky130_fd_sc_hd__or2b_1
X_12385_ net572 _05230_ _05233_ _05234_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14124_ _06836_ _06838_ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_244_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19981_ _01563_ _01780_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14055_ top_inst.grid_inst.data_path_wires\[3\]\[0\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _06771_ sky130_fd_sc_hd__or2b_1
XFILLER_0_162_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18932_ _11164_ _11132_ _11316_ VGND VGND VPWR VPWR _11355_ sky130_fd_sc_hd__and3_1
XFILLER_0_205_1388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13006_ top_inst.grid_inst.data_path_wires\[1\]\[1\] top_inst.grid_inst.data_path_wires\[1\]\[0\]
+ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[3\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[2\]
+ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18863_ _11258_ _11259_ _11286_ _11287_ VGND VGND VPWR VPWR _11288_ sky130_fd_sc_hd__a211o_1
XTAP_6560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17814_ _10278_ _10320_ _09292_ VGND VGND VPWR VPWR _10322_ sky130_fd_sc_hd__a21o_1
XTAP_6593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18794_ _11217_ _11220_ VGND VGND VPWR VPWR _11221_ sky130_fd_sc_hd__xor2_2
XFILLER_0_94_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17745_ _10244_ _10253_ VGND VGND VPWR VPWR _10254_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_206_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14957_ _04865_ _07460_ VGND VGND VPWR VPWR _07623_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13908_ _05260_ VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__clkbuf_4
X_17676_ _10184_ _10185_ _10147_ _10146_ VGND VGND VPWR VPWR _10187_ sky130_fd_sc_hd__o2bb2a_1
X_14888_ _07570_ _07571_ VGND VGND VPWR VPWR _07572_ sky130_fd_sc_hd__and2_1
XFILLER_0_187_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19415_ _01247_ _01248_ _01249_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__o21bai_2
X_16627_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _09198_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13839_ _06548_ _06551_ _06580_ VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__and3_1
XFILLER_0_230_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_230_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19346_ _11693_ _11677_ _11682_ _11688_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16558_ _09116_ _09099_ _09132_ VGND VGND VPWR VPWR _09134_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15509_ _07613_ _06634_ _08144_ _08142_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19277_ _09185_ _11677_ _11680_ _11641_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16489_ _09028_ _09030_ VGND VGND VPWR VPWR _09067_ sky130_fd_sc_hd__or2b_1
XFILLER_0_127_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18228_ _10692_ _10696_ VGND VGND VPWR VPWR _10697_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18159_ _10629_ _10630_ VGND VGND VPWR VPWR _10631_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold302 _00213_ VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold313 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[0\] VGND
+ VGND VPWR VPWR net495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[29\] VGND
+ VGND VPWR VPWR net506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 top_inst.axis_out_inst.out_buff_data\[118\] VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21170_ _02911_ _02912_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__nand2_1
Xhold346 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[7\] VGND
+ VGND VPWR VPWR net528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 _00149_ VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20121_ _01916_ _01920_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__nand2_1
Xhold368 _00084_ VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold379 top_inst.deskew_buff_inst.col_input\[93\] VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_141_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20052_ _01824_ _01866_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23811_ clknet_leaf_72_clk _00344_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_240_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23742_ clknet_leaf_127_clk net450 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20954_ _02688_ _02722_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23673_ clknet_leaf_116_clk _00206_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_20885_ _02624_ _02642_ _02655_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__nand3_1
XFILLER_0_49_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_634 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22624_ _04299_ _04300_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__and2_1
XFILLER_0_187_1314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22555_ _04208_ _04211_ _04234_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21506_ _03227_ _03229_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22486_ _04166_ _04167_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24225_ clknet_leaf_112_clk _00758_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[16\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21437_ _02873_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[5\] VGND
+ VGND VPWR VPWR _03172_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24156_ clknet_leaf_17_clk _00689_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12170_ net566 _05110_ _05111_ _05101_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__o211a_1
X_21368_ _03074_ _03104_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__xor2_2
XFILLER_0_20_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23107_ top_inst.valid_pipe\[7\] _05323_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20319_ top_inst.grid_inst.data_path_wires\[16\]\[5\] _01986_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[5\]
+ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _02107_ sky130_fd_sc_hd__and4_1
XFILLER_0_198_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24087_ clknet_leaf_86_clk _00620_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold880 top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[14\] VGND VGND
+ VPWR VPWR net1062 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21299_ _03012_ _03013_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__nor2_1
Xhold891 top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[3\] VGND VGND
+ VPWR VPWR net1073 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23038_ top_inst.axis_in_inst.inbuf_bus\[9\] _04603_ VGND VGND VPWR VPWR _04614_
+ sky130_fd_sc_hd__or2_1
XTAP_5100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15860_ _08469_ _08471_ _08265_ VGND VGND VPWR VPWR _08473_ sky130_fd_sc_hd__o21a_1
XFILLER_0_244_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14811_ _07241_ _07085_ _07496_ VGND VGND VPWR VPWR _07497_ sky130_fd_sc_hd__or3_1
XTAP_5188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _08147_ _08164_ _08161_ _08149_ VGND VGND VPWR VPWR _08405_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _10029_ _10046_ _10051_ _10049_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__o211a_1
X_14742_ _07387_ _07389_ VGND VGND VPWR VPWR _07430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11954_ net699 _04982_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_1112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14673_ _07349_ _07318_ VGND VGND VPWR VPWR _07362_ sky130_fd_sc_hd__or2b_4
X_17461_ _09995_ _09996_ VGND VGND VPWR VPWR _09997_ sky130_fd_sc_hd__and2_1
XFILLER_0_200_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11885_ net800 _04943_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__or2_1
XFILLER_0_170_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19200_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[14\] _10639_ VGND
+ VGND VPWR VPWR _11617_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16412_ _08990_ _08991_ VGND VGND VPWR VPWR _08992_ sky130_fd_sc_hd__nor2_1
X_13624_ _06369_ _06370_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17392_ _09910_ _09908_ _09925_ VGND VGND VPWR VPWR _09931_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_131_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19131_ _11506_ _11507_ _11539_ VGND VGND VPWR VPWR _11549_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16343_ _08695_ _08671_ VGND VGND VPWR VPWR _08924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13555_ _06294_ _06303_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_229_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12506_ top_inst.axis_in_inst.inbuf_valid _05323_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__nand2_1
X_16274_ _08855_ _08856_ VGND VGND VPWR VPWR _08857_ sky130_fd_sc_hd__xnor2_1
X_19062_ _11480_ _11481_ _11145_ _11161_ VGND VGND VPWR VPWR _11482_ sky130_fd_sc_hd__and4b_1
XFILLER_0_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13486_ _06186_ _06217_ _06219_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__nor3_1
XFILLER_0_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15225_ _07870_ _07871_ VGND VGND VPWR VPWR _07872_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18013_ _10479_ _10515_ VGND VGND VPWR VPWR _10516_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_180_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12437_ net300 _05256_ _05264_ _05261_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15156_ _07803_ _07804_ VGND VGND VPWR VPWR _07805_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12368_ net835 _05222_ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14107_ _06741_ _06774_ _06821_ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19964_ _01611_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__clkbuf_4
X_15087_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[5\] _06242_ _07736_
+ _07737_ VGND VGND VPWR VPWR _07738_ sky130_fd_sc_hd__a22o_1
X_12299_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[4\] _05183_
+ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__or2_1
XFILLER_0_226_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14038_ _06717_ _06754_ VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__xnor2_2
X_18915_ _11152_ _11149_ _11147_ VGND VGND VPWR VPWR _11338_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_238_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19895_ _01715_ _01711_ _01716_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18846_ _11231_ _11236_ VGND VGND VPWR VPWR _11271_ sky130_fd_sc_hd__or2b_1
XTAP_6390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18777_ _11190_ _11203_ _11204_ VGND VGND VPWR VPWR _11205_ sky130_fd_sc_hd__nand3_1
XFILLER_0_171_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15989_ _08595_ _08596_ _08517_ _08597_ VGND VGND VPWR VPWR _08598_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_171_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17728_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[8\] _10236_ VGND
+ VGND VPWR VPWR _10237_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17659_ _10168_ _10169_ VGND VGND VPWR VPWR _10170_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20670_ _02447_ _02449_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__xor2_1
XFILLER_0_174_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19329_ _05326_ VGND VGND VPWR VPWR _11723_ sky130_fd_sc_hd__buf_6
XFILLER_0_45_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22340_ _03693_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[5\] VGND
+ VGND VPWR VPWR _04026_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22271_ _03956_ _03958_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__xor2_2
XFILLER_0_108_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24010_ clknet_leaf_47_clk _00543_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold110 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[20\] VGND
+ VGND VPWR VPWR net292 sky130_fd_sc_hd__dlygate4sd3_1
X_21222_ net604 _02491_ _02960_ _02961_ _02962_ VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__o221a_1
Xhold121 _01159_ VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold132 _00042_ VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 top_inst.deskew_buff_inst.col_input\[65\] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _00293_ VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _00183_ VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__dlygate4sd3_1
X_21153_ _02878_ _02881_ _02898_ _02880_ VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__o211a_1
Xhold176 _00177_ VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[27\] VGND
+ VGND VPWR VPWR net369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold198 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[6\] VGND VGND
+ VPWR VPWR net380 sky130_fd_sc_hd__dlygate4sd3_1
X_20104_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[28\] _01764_ VGND
+ VGND VPWR VPWR _01917_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_217_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21084_ _02845_ _02846_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20035_ _01783_ _01831_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21986_ top_inst.grid_inst.data_path_wires\[18\]\[6\] VGND VGND VPWR VPWR _03693_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_240_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23725_ clknet_leaf_136_clk net307 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20937_ _02706_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23656_ clknet_leaf_132_clk net353 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20868_ _02614_ _02631_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_667 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22607_ _04188_ _04254_ _04281_ _04282_ _04283_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_181_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23587_ clknet_leaf_105_clk net281 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20799_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[18\] _02467_ VGND
+ VGND VPWR VPWR _02574_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13340_ _06095_ _06099_ _06093_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__o21a_1
XFILLER_0_221_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22538_ _04061_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__buf_2
XFILLER_0_10_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13271_ _05751_ _05768_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__nand2_1
XFILLER_0_224_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22469_ _04118_ _04151_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__xor2_1
XFILLER_0_49_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15010_ _07662_ _07663_ VGND VGND VPWR VPWR _07664_ sky130_fd_sc_hd__and2_1
X_24208_ clknet_leaf_17_clk _00741_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12222_ net343 _05137_ _05140_ _05141_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__o211a_1
XFILLER_0_224_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12153_ _05009_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__buf_2
X_24139_ clknet_leaf_4_clk _00672_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[25\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_103_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16961_ _09513_ net220 _09515_ VGND VGND VPWR VPWR _09516_ sky130_fd_sc_hd__nand3_1
X_12084_ _05009_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_159_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_235_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18700_ _10583_ VGND VGND VPWR VPWR _11142_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15912_ _08150_ _08167_ _08486_ _08485_ VGND VGND VPWR VPWR _08523_ sky130_fd_sc_hd__a31o_1
X_19680_ _01508_ _01509_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__xnor2_2
X_16892_ _09447_ _09448_ VGND VGND VPWR VPWR _09449_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_232_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18631_ _11088_ _11089_ VGND VGND VPWR VPWR _11090_ sky130_fd_sc_hd__or2_1
XTAP_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ _08454_ _08455_ VGND VGND VPWR VPWR _08456_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_239_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_235_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18562_ _11021_ _11022_ VGND VGND VPWR VPWR _11023_ sky130_fd_sc_hd__nand2_1
XTAP_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[7\] _05773_ VGND
+ VGND VPWR VPWR _05774_ sky130_fd_sc_hd__or2_1
XTAP_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ _08333_ _08334_ _08388_ VGND VGND VPWR VPWR _08389_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17513_ _10038_ _10033_ _10039_ _10024_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__o211a_1
X_14725_ _07079_ _07074_ _07090_ VGND VGND VPWR VPWR _07413_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_185_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ net520 _04977_ _04978_ _04968_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__o211a_1
X_18493_ _10914_ _10917_ _10955_ VGND VGND VPWR VPWR _10956_ sky130_fd_sc_hd__a21oi_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _09919_ _09957_ _09937_ VGND VGND VPWR VPWR _09981_ sky130_fd_sc_hd__or3b_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14656_ _07344_ _07345_ VGND VGND VPWR VPWR _07346_ sky130_fd_sc_hd__and2_2
XFILLER_0_157_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11868_ net753 _04938_ _04939_ _04929_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13607_ _06353_ _06354_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__xnor2_1
X_17375_ _09913_ _09914_ VGND VGND VPWR VPWR _09915_ sky130_fd_sc_hd__nand2_2
XFILLER_0_7_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14587_ _07066_ _07062_ _07090_ VGND VGND VPWR VPWR _07278_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_32_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11799_ top_inst.axis_out_inst.out_buff_data\[78\] _04890_ VGND VGND VPWR VPWR _04900_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_55_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19114_ _11479_ _11487_ _11532_ VGND VGND VPWR VPWR _11533_ sky130_fd_sc_hd__a21bo_1
X_16326_ _08905_ _08907_ VGND VGND VPWR VPWR _08908_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13538_ _05886_ _06287_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19045_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[10\] _10639_ VGND
+ VGND VPWR VPWR _11466_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16257_ _08693_ top_inst.grid_inst.data_path_wires\[8\]\[4\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[3\]
+ _08669_ VGND VGND VPWR VPWR _08840_ sky130_fd_sc_hd__nand4_2
X_13469_ net1004 _05788_ _06222_ _06207_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15208_ _07853_ _07855_ VGND VGND VPWR VPWR _07856_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16188_ top_inst.grid_inst.data_path_wires\[8\]\[4\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[1\]
+ _08682_ top_inst.grid_inst.data_path_wires\[8\]\[5\] VGND VGND VPWR VPWR _08773_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_199_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15139_ top_inst.grid_inst.data_path_wires\[6\]\[4\] top_inst.grid_inst.data_path_wires\[6\]\[3\]
+ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _07788_ sky130_fd_sc_hd__nand4_2
XFILLER_0_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19947_ _01561_ _01765_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19878_ _01698_ _01700_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_177_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_896 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18829_ _11229_ _11253_ _10831_ VGND VGND VPWR VPWR _11255_ sky130_fd_sc_hd__o21a_1
XFILLER_0_223_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21840_ _03560_ _03551_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_223_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21771_ _03493_ _03494_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23510_ clknet_leaf_137_clk _00043_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20722_ _02498_ _02499_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24490_ clknet_leaf_45_clk _01023_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_enabled
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23441_ net659 _04840_ _04842_ _04831_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20653_ _02001_ _02229_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23372_ _04686_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__buf_2
XFILLER_0_11_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20584_ _02364_ _02365_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_85_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22323_ top_inst.deskew_buff_inst.col_input\[106\] _05731_ _04008_ _04009_ VGND VGND
+ VPWR VPWR _04010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22254_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[9\] _03894_ VGND
+ VGND VPWR VPWR _03942_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21205_ _02944_ _02945_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__nand2_1
X_22185_ _03849_ _03874_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__xor2_1
XFILLER_0_160_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21136_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _02887_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_217_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21067_ _02503_ _02793_ _02812_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__or3_1
X_20018_ _01809_ _01833_ _01826_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__nand3_1
XFILLER_0_236_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12840_ _05645_ _05646_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__nor2_1
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_241_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _05564_ _05540_ _05578_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__nand3_1
XFILLER_0_198_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21969_ _02862_ _02877_ _03681_ _03660_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__o211a_1
XFILLER_0_240_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[2\] _07078_ _07200_
+ _07201_ VGND VGND VPWR VPWR _07203_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_1126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15490_ _08126_ _08129_ VGND VGND VPWR VPWR _08130_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23708_ clknet_leaf_124_clk _00241_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[1\] _07072_ _07077_
+ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _07136_ sky130_fd_sc_hd__a22o_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23639_ clknet_leaf_126_clk _00172_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14372_ _07074_ _07075_ VGND VGND VPWR VPWR _07076_ sky130_fd_sc_hd__or2_1
X_17160_ _09707_ _09709_ VGND VGND VPWR VPWR _09710_ sky130_fd_sc_hd__xor2_1
XFILLER_0_154_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13323_ _06096_ _06016_ net182 VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__or3_2
X_16111_ _08683_ _08661_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _08701_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17091_ _09640_ _09641_ _09553_ VGND VGND VPWR VPWR _09643_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_162_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13254_ _06028_ _06030_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__xor2_1
XFILLER_0_122_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16042_ _08627_ _08635_ VGND VGND VPWR VPWR _08649_ sky130_fd_sc_hd__or2_1
XFILLER_0_204_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12205_ top_inst.axis_out_inst.out_buff_data\[28\] _05129_ VGND VGND VPWR VPWR _05132_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_122_1109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13185_ _05925_ _05921_ _05962_ _05405_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_86_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19801_ _01626_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__inv_2
XFILLER_0_236_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12136_ net823 _05084_ _05092_ _05088_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17993_ _10490_ _10494_ VGND VGND VPWR VPWR _10496_ sky130_fd_sc_hd__or2_1
XFILLER_0_202_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19732_ _01552_ _01520_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__or2b_1
X_16944_ _09460_ _09463_ _09498_ VGND VGND VPWR VPWR _09499_ sky130_fd_sc_hd__a21o_1
X_12067_ net877 _05045_ _05053_ _05049_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__o211a_1
X_19663_ _01490_ _01491_ _01489_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__a21o_1
X_16875_ _09429_ _09430_ _09428_ VGND VGND VPWR VPWR _09432_ sky130_fd_sc_hd__a21o_1
XFILLER_0_204_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18614_ _11033_ _11069_ VGND VGND VPWR VPWR _11073_ sky130_fd_sc_hd__or2b_1
XTAP_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15826_ _08437_ _08438_ VGND VGND VPWR VPWR _08439_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19594_ _01424_ _01425_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__and2_1
XTAP_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18545_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[12\] _10923_ _10840_
+ VGND VGND VPWR VPWR _11006_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_138_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_138_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15757_ top_inst.grid_inst.data_path_wires\[7\]\[7\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _08372_ sky130_fd_sc_hd__and3_1
XTAP_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _05761_ _05294_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__or2_1
XTAP_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14708_ _07394_ _07395_ _07361_ _07362_ VGND VGND VPWR VPWR _07397_ sky130_fd_sc_hd__o211a_1
X_18476_ _10936_ _10938_ VGND VGND VPWR VPWR _10939_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15688_ _08211_ _08233_ _08260_ _08264_ VGND VGND VPWR VPWR _08305_ sky130_fd_sc_hd__o31a_1
XFILLER_0_157_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17427_ _09963_ _09964_ VGND VGND VPWR VPWR _09965_ sky130_fd_sc_hd__nor2_1
X_14639_ _07079_ _07082_ _07086_ _07074_ VGND VGND VPWR VPWR _07329_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17358_ _09894_ _09898_ VGND VGND VPWR VPWR _09899_ sky130_fd_sc_hd__xor2_2
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16309_ _08798_ _08837_ _08890_ VGND VGND VPWR VPWR _08891_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_127_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17289_ _09813_ _09815_ _09832_ VGND VGND VPWR VPWR _09833_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19028_ _11441_ _11448_ VGND VGND VPWR VPWR _11449_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23990_ clknet_leaf_78_clk _00523_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_103_1097 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22941_ net1015 _04548_ _04558_ _04551_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_1116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22872_ top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[2\] _04517_ VGND
+ VGND VPWR VPWR _04519_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24611_ clknet_leaf_21_clk _01144_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_151_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21823_ net670 _03528_ _03543_ _03544_ _02962_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__o221a_1
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_129_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_129_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_222_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24542_ clknet_leaf_100_clk _01075_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dfxtp_4
X_21754_ _03478_ _03470_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20705_ _02425_ _02445_ _02444_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__o21ba_1
X_24473_ clknet_leaf_37_clk _01006_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21685_ _03372_ _03386_ _03384_ VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_188_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_946 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23424_ top_inst.axis_out_inst.out_buff_data\[101\] _04596_ VGND VGND VPWR VPWR _04833_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_135_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20636_ _02391_ _02392_ _02415_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__nand3_1
XFILLER_0_164_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_862 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23355_ net41 _04792_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20567_ _02349_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22306_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[5\] _03688_ _03955_
+ _03992_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23286_ net135 _04753_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__or2_1
X_20498_ _02274_ _02281_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__xor2_1
XFILLER_0_225_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22237_ _03923_ _03925_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__xor2_2
XFILLER_0_218_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22168_ _03850_ _03856_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__or2_1
XFILLER_0_218_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21119_ _01999_ _11142_ _02874_ _02707_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__o211a_1
XFILLER_0_234_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14990_ _07606_ _07627_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _07646_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22099_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[5\] _03790_ VGND
+ VGND VPWR VPWR _03791_ sky130_fd_sc_hd__xor2_2
XFILLER_0_233_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13941_ _06656_ _06661_ VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__or2_1
XFILLER_0_233_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_242_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16660_ _09194_ _09187_ _09192_ _09189_ VGND VGND VPWR VPWR _09224_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13872_ _06555_ _06599_ _06597_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_214_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_236_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15611_ _08225_ _08229_ VGND VGND VPWR VPWR _08230_ sky130_fd_sc_hd__xor2_2
X_12823_ _05629_ _05630_ _05328_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__a21o_1
XFILLER_0_243_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16591_ _09163_ _09164_ VGND VGND VPWR VPWR _09166_ sky130_fd_sc_hd__and2_1
XFILLER_0_201_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_863 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18330_ _10789_ _10795_ VGND VGND VPWR VPWR _10796_ sky130_fd_sc_hd__xnor2_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15542_ _08167_ _07641_ VGND VGND VPWR VPWR _08168_ sky130_fd_sc_hd__or2_1
X_12754_ _05542_ _05544_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18261_ top_inst.grid_inst.data_path_wires\[12\]\[3\] top_inst.grid_inst.data_path_wires\[12\]\[2\]
+ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _10729_ sky130_fd_sc_hd__and4_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _05494_ _05495_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__xnor2_2
X_15473_ _08112_ _08113_ VGND VGND VPWR VPWR _08114_ sky130_fd_sc_hd__or2_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17212_ _09751_ _09759_ VGND VGND VPWR VPWR _09760_ sky130_fd_sc_hd__xor2_1
X_14424_ _07066_ _07062_ _07069_ _07073_ VGND VGND VPWR VPWR _07120_ sky130_fd_sc_hd__nand4_1
XFILLER_0_182_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18192_ _10641_ _10662_ VGND VGND VPWR VPWR _10663_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17143_ _09691_ _09693_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[14\]
+ _07816_ VGND VGND VPWR VPWR _09694_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_167_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14355_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _07062_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13306_ _06049_ _06048_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__or2b_1
X_17074_ _09625_ _09592_ VGND VGND VPWR VPWR _09626_ sky130_fd_sc_hd__nor2_1
X_14286_ _06976_ _06980_ _06974_ VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__o21a_1
Xhold709 top_inst.deskew_buff_inst.col_input\[81\] VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13237_ _05970_ _05973_ _05971_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_21_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16025_ _08628_ _08632_ VGND VGND VPWR VPWR _08633_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13168_ _05896_ _05898_ _05946_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_1340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12119_ net264 _05071_ _05082_ _05075_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__o211a_1
XFILLER_0_237_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13099_ _05874_ _05875_ _05878_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__o21a_1
X_17976_ _10477_ _10478_ VGND VGND VPWR VPWR _10480_ sky130_fd_sc_hd__nand2_1
XFILLER_0_236_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19715_ _01541_ _01542_ _01543_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__nand3_1
XFILLER_0_139_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16927_ net200 _09481_ _09482_ VGND VGND VPWR VPWR _09483_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19646_ _01436_ _01439_ _01475_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__a21o_1
X_16858_ _09198_ _09210_ _09374_ _09373_ VGND VGND VPWR VPWR _09415_ sky130_fd_sc_hd__a31o_1
XFILLER_0_215_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15809_ _08369_ _08381_ _08422_ VGND VGND VPWR VPWR _08423_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_1062 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19577_ _01298_ _11686_ net239 _11703_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_137_1182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16789_ _09300_ _09302_ _09346_ _09347_ VGND VGND VPWR VPWR _09348_ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18528_ _10974_ _10989_ VGND VGND VPWR VPWR _10990_ sky130_fd_sc_hd__xor2_1
XFILLER_0_158_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_220_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18459_ _10885_ _10888_ _10921_ VGND VGND VPWR VPWR _10922_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_185_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21470_ _03202_ _03203_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20421_ _02204_ _02205_ _02160_ _02162_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23140_ net49 _04672_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__or2_1
X_20352_ _02107_ _02137_ _02138_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__and3_1
XFILLER_0_222_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23071_ net15 _04628_ _04633_ _04632_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__o211a_1
X_20283_ _05312_ _02070_ _02071_ _02072_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22022_ _03682_ _03698_ _03680_ _03700_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__a22o_1
XTAP_6219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23973_ clknet_leaf_86_clk _00506_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_231_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22924_ _10583_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_230_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22855_ _10583_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_210_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21806_ _06168_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22786_ _04192_ _04412_ _04431_ _04434_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__a31o_1
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24525_ clknet_leaf_128_clk _01058_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dfxtp_4
X_21737_ _03433_ _03462_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12470_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _05293_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24456_ clknet_4_15__leaf_clk _00989_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21668_ _03341_ _03395_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23407_ net67 _04658_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20619_ _01999_ _02229_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__nor2_1
X_24387_ clknet_leaf_38_clk net388 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21599_ _03210_ _03329_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__xnor2_2
X_14140_ _06852_ _06853_ VGND VGND VPWR VPWR _06854_ sky130_fd_sc_hd__xnor2_1
X_23338_ net160 _04779_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_1362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14071_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[7\] _06784_ _06786_
+ VGND VGND VPWR VPWR _06787_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23269_ net127 _04740_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13022_ top_inst.grid_inst.data_path_wires\[1\]\[3\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[1\]\[4\]
+ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__a22o_1
XTAP_6720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17830_ _10038_ _10335_ _10336_ VGND VGND VPWR VPWR _10337_ sky130_fd_sc_hd__a21bo_1
XTAP_6753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17761_ _10266_ _10268_ VGND VGND VPWR VPWR _10270_ sky130_fd_sc_hd__and2_1
X_14973_ _07633_ _07075_ VGND VGND VPWR VPWR _07634_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19500_ _01330_ _01331_ _01332_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__o21ai_2
X_16712_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[3\] _09248_ _09249_
+ VGND VGND VPWR VPWR _09273_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_57_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13924_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _06650_ sky130_fd_sc_hd__clkbuf_4
X_17692_ _10197_ _10201_ VGND VGND VPWR VPWR _10202_ sky130_fd_sc_hd__xor2_2
XFILLER_0_107_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19431_ _01239_ _01240_ _01264_ _01265_ VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__a211o_1
X_16643_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _09211_ sky130_fd_sc_hd__buf_2
XFILLER_0_186_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13855_ _06541_ _06595_ VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12806_ _05611_ _05613_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19362_ _05887_ _01197_ _01198_ _01199_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16574_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[15\] _05634_ VGND
+ VGND VPWR VPWR _09149_ sky130_fd_sc_hd__and2_1
XFILLER_0_202_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13786_ _06525_ _06526_ VGND VGND VPWR VPWR _06529_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18313_ _10614_ _10779_ VGND VGND VPWR VPWR _10780_ sky130_fd_sc_hd__xnor2_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15525_ _08155_ _07641_ VGND VGND VPWR VPWR _08156_ sky130_fd_sc_hd__or2_1
X_12737_ _05507_ _05546_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__or2_1
X_19293_ _11693_ _11689_ VGND VGND VPWR VPWR _11694_ sky130_fd_sc_hd__or2_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18244_ _10700_ _10702_ VGND VGND VPWR VPWR _10712_ sky130_fd_sc_hd__nand2_1
X_15456_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[14\] _08066_ _08096_
+ _08097_ VGND VGND VPWR VPWR _08098_ sky130_fd_sc_hd__a22o_1
X_12668_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[7\] _05326_ VGND
+ VGND VPWR VPWR _05480_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14407_ _07066_ _07062_ _07065_ _07069_ VGND VGND VPWR VPWR _07104_ sky130_fd_sc_hd__nand4_2
X_18175_ _10602_ _10645_ VGND VGND VPWR VPWR _10646_ sky130_fd_sc_hd__nand2_2
X_15387_ _07995_ _07996_ VGND VGND VPWR VPWR _08030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12599_ _05377_ _05382_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17126_ _09551_ _09552_ _09674_ _09675_ VGND VGND VPWR VPWR _09677_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_106_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14338_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[14\] _05634_ _07045_
+ _07046_ VGND VGND VPWR VPWR _07047_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold506 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[27\] VGND
+ VGND VPWR VPWR net688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold517 top_inst.axis_out_inst.out_buff_data\[49\] VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold528 top_inst.axis_out_inst.out_buff_data\[112\] VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__dlygate4sd3_1
X_17057_ _09607_ _09608_ _09594_ VGND VGND VPWR VPWR _09610_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold539 _00098_ VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__dlygate4sd3_1
X_14269_ _06978_ _06979_ VGND VGND VPWR VPWR _06980_ sky130_fd_sc_hd__nand2_2
XFILLER_0_141_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16008_ _08614_ _08616_ VGND VGND VPWR VPWR _08617_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ _10419_ _10462_ VGND VGND VPWR VPWR _10463_ sky130_fd_sc_hd__xnor2_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20970_ net696 _02638_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__or2_1
XFILLER_0_212_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19629_ _01418_ _01435_ _01458_ _01459_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__a211o_1
XFILLER_0_221_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22640_ _04306_ _04314_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22571_ _04248_ _04249_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__and2_1
XFILLER_0_186_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24310_ clknet_leaf_2_clk _00843_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[85\]
+ sky130_fd_sc_hd__dfxtp_1
X_21522_ top_inst.grid_inst.data_path_wires\[17\]\[6\] _02895_ VGND VGND VPWR VPWR
+ _03255_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_1036 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24241_ clknet_leaf_112_clk _00774_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21453_ _03162_ _03187_ VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20404_ _01992_ _02018_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24172_ clknet_leaf_23_clk _00705_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21384_ _03075_ _03082_ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23123_ net677 _04656_ _04663_ _04662_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20335_ _02104_ _02105_ _02120_ _02121_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_113_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1081 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput37 net37 VGND VGND VPWR VPWR input_tready sky130_fd_sc_hd__clkbuf_4
XTAP_6005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23054_ net7 _04615_ _04623_ _04619_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__o211a_1
X_20266_ _02038_ _02054_ _02055_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__or3b_2
Xoutput48 net48 VGND VGND VPWR VPWR output_tdata[109] sky130_fd_sc_hd__clkbuf_4
Xoutput59 net59 VGND VGND VPWR VPWR output_tdata[119] sky130_fd_sc_hd__clkbuf_4
XTAP_6016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22005_ _03686_ _05270_ _03706_ _03702_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__o211a_1
XTAP_6049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20197_ _01999_ _10033_ _02000_ _01840_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__o211a_1
XTAP_5337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23956_ clknet_leaf_91_clk _00489_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11970_ top_inst.axis_out_inst.out_buff_data\[55\] _04996_ VGND VGND VPWR VPWR _04998_
+ sky130_fd_sc_hd__or2_1
XTAP_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22907_ top_inst.skew_buff_inst.row\[2\].output_reg\[1\] _04530_ VGND VGND VPWR VPWR
+ _04539_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23887_ clknet_leaf_64_clk _00420_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13640_ _06335_ _06337_ _06386_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__a21o_1
X_22838_ top_inst.skew_buff_inst.row\[3\].output_reg\[3\] _03691_ VGND VGND VPWR VPWR
+ _04500_ sky130_fd_sc_hd__or2_1
XFILLER_0_233_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_838 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ _06315_ _06316_ _06319_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__nor3_2
XFILLER_0_183_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22769_ _04436_ _04437_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__and2_1
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_51_clk clknet_4_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15310_ _07916_ _07954_ VGND VGND VPWR VPWR _07955_ sky130_fd_sc_hd__nor2_2
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12522_ _05288_ _05272_ _05279_ _05284_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_13_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24508_ clknet_leaf_127_clk _01041_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dfxtp_4
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16290_ _08864_ _08865_ _08871_ VGND VGND VPWR VPWR _08872_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15241_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[9\] _07845_ VGND
+ VGND VPWR VPWR _07888_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24439_ clknet_leaf_58_clk net584 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12453_ _05278_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15172_ _07812_ _07813_ _07819_ VGND VGND VPWR VPWR _07820_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12384_ _05127_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__buf_2
XFILLER_0_65_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_240_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14123_ _06751_ _06790_ _06837_ VGND VGND VPWR VPWR _06838_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_22_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19980_ _01792_ _01795_ net168 VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18931_ _11349_ _11353_ VGND VGND VPWR VPWR _11354_ sky130_fd_sc_hd__xnor2_1
X_14054_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[3\]\[1\]
+ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__nand2_1
XFILLER_0_219_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13005_ _05734_ _05763_ _05761_ _05738_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_120_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18862_ _11284_ _11285_ _11260_ _11261_ VGND VGND VPWR VPWR _11287_ sky130_fd_sc_hd__o211a_1
XTAP_6550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17813_ _10278_ _10320_ VGND VGND VPWR VPWR _10321_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18793_ _11218_ _11219_ VGND VGND VPWR VPWR _11220_ sky130_fd_sc_hd__nand2_1
XTAP_5860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17744_ _10250_ _10252_ VGND VGND VPWR VPWR _10253_ sky130_fd_sc_hd__xnor2_1
XTAP_5893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14956_ _07621_ VGND VGND VPWR VPWR _07622_ sky130_fd_sc_hd__buf_4
XFILLER_0_221_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13907_ _06637_ _05773_ VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__or2_1
XFILLER_0_216_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17675_ _10147_ _10146_ _10184_ _10185_ VGND VGND VPWR VPWR _10186_ sky130_fd_sc_hd__and4bb_1
X_14887_ _07540_ _07544_ _07569_ VGND VGND VPWR VPWR _07571_ sky130_fd_sc_hd__nand3_1
XFILLER_0_221_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19414_ _01247_ _01248_ _01249_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__or3b_4
X_16626_ net224 VGND VGND VPWR VPWR _09197_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_173_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13838_ _06578_ _06579_ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__nand2_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19345_ _11724_ _11731_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16557_ _09116_ _09099_ _09132_ VGND VGND VPWR VPWR _09133_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13769_ _06510_ _06511_ VGND VGND VPWR VPWR _06513_ sky130_fd_sc_hd__and2_1
XFILLER_0_186_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_42_clk clknet_4_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15508_ _08143_ _08140_ VGND VGND VPWR VPWR _08144_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19276_ _11679_ _11150_ VGND VGND VPWR VPWR _11680_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16488_ _09063_ _09065_ VGND VGND VPWR VPWR _09066_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18227_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[5\] _10695_ VGND
+ VGND VPWR VPWR _10696_ sky130_fd_sc_hd__xor2_2
X_15439_ _08079_ _08080_ VGND VGND VPWR VPWR _08081_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18158_ _10581_ _10599_ _10600_ _10597_ VGND VGND VPWR VPWR _10630_ sky130_fd_sc_hd__nand4_1
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold303 top_inst.axis_out_inst.out_buff_data\[17\] VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17109_ net1049 _09266_ _09659_ _09660_ _07708_ VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__o221a_1
XFILLER_0_124_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold314 _00263_ VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold325 _00164_ VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__dlygate4sd3_1
X_18089_ _10022_ _08663_ _10578_ _10448_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold336 top_inst.deskew_buff_inst.col_input\[63\] VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__buf_1
XFILLER_0_1_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold347 _00238_ VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20120_ _01912_ _01929_ _01927_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__a21boi_1
Xhold358 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[21\] VGND
+ VGND VPWR VPWR net540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold369 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[28\] VGND
+ VGND VPWR VPWR net551 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_3__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_4_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_229_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20051_ _01865_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__inv_2
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23810_ clknet_leaf_72_clk _00343_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20953_ _02720_ _02721_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__nor2_1
X_23741_ clknet_leaf_122_clk net536 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ _02624_ _02642_ _02655_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__a21o_1
X_23672_ clknet_leaf_116_clk _00205_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22623_ _04275_ _04298_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__or2_1
XFILLER_0_193_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_33_clk clknet_4_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_187_1326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22554_ _04205_ _04233_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__xor2_1
XFILLER_0_174_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21505_ _03191_ _03235_ _03236_ _03072_ _03237_ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_161_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22485_ _04061_ _04165_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24224_ clknet_leaf_19_clk _00757_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21436_ _03135_ _03170_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__xor2_2
XFILLER_0_133_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24155_ clknet_leaf_18_clk _00688_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21367_ _03101_ _03103_ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23106_ net354 _10541_ _04651_ _04643_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__o211a_1
X_20318_ _01987_ _02018_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[0\]
+ _01999_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__a22oi_1
X_24086_ clknet_leaf_87_clk _00619_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold870 top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[11\] VGND VGND
+ VPWR VPWR net1052 sky130_fd_sc_hd__dlygate4sd3_1
X_21298_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[6\] _03000_ _03001_
+ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__a21bo_1
Xhold881 top_inst.skew_buff_inst.row\[0\].output_reg\[6\] VGND VGND VPWR VPWR net1063
+ sky130_fd_sc_hd__dlygate4sd3_1
X_23037_ net31 _04601_ _04613_ _04606_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold892 top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[15\] VGND VGND
+ VPWR VPWR net1074 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20249_ _02037_ _02038_ _02039_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_219_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _07087_ _07089_ VGND VGND VPWR VPWR _07496_ sky130_fd_sc_hd__nand2_1
XTAP_5178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _08402_ _08403_ VGND VGND VPWR VPWR _08404_ sky130_fd_sc_hd__xor2_1
XTAP_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14741_ _07409_ _07427_ VGND VGND VPWR VPWR _07429_ sky130_fd_sc_hd__nand2_1
XTAP_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23939_ clknet_leaf_81_clk _00472_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ net967 _04977_ _04987_ _04981_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__o211a_1
XTAP_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17460_ _09913_ _09974_ _09994_ VGND VGND VPWR VPWR _09996_ sky130_fd_sc_hd__nand3_1
XTAP_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _07346_ _07348_ VGND VGND VPWR VPWR _07361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_1352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11884_ net503 _04938_ _04948_ _04942_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__o211a_1
XFILLER_0_197_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16411_ _08952_ _08989_ VGND VGND VPWR VPWR _08991_ sky130_fd_sc_hd__nor2_1
XFILLER_0_200_956 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_184_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13623_ _06188_ _06212_ VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17391_ _09929_ VGND VGND VPWR VPWR _09930_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_clk clknet_4_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19130_ _11498_ _11540_ _11541_ VGND VGND VPWR VPWR _11548_ sky130_fd_sc_hd__or3_1
X_16342_ _08921_ _08922_ VGND VGND VPWR VPWR _08923_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13554_ _06297_ _06302_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19061_ _11351_ _11140_ _11143_ _11164_ VGND VGND VPWR VPWR _11481_ sky130_fd_sc_hd__a2bb2o_1
X_12505_ _05267_ _04856_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__nor2_2
XFILLER_0_192_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16273_ _08796_ _08805_ _08815_ VGND VGND VPWR VPWR _08856_ sky130_fd_sc_hd__o21ai_1
X_13485_ _06231_ _06236_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18012_ _10511_ _10514_ VGND VGND VPWR VPWR _10515_ sky130_fd_sc_hd__xor2_2
X_15224_ top_inst.grid_inst.data_path_wires\[6\]\[3\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[6\]
+ _07824_ top_inst.grid_inst.data_path_wires\[6\]\[2\] VGND VGND VPWR VPWR _07871_
+ sky130_fd_sc_hd__o2bb2a_1
X_12436_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[31\] _05262_
+ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__or2_1
XFILLER_0_242_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15155_ _07717_ _07753_ _07764_ VGND VGND VPWR VPWR _07804_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12367_ net466 _05217_ _05224_ _05221_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14106_ _06775_ _06778_ _06779_ VGND VGND VPWR VPWR _06821_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19963_ _01779_ _01781_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__xor2_2
X_15086_ _07709_ _07735_ _05315_ VGND VGND VPWR VPWR _07737_ sky130_fd_sc_hd__o21a_1
X_12298_ net494 _05178_ _05185_ _05182_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14037_ _06750_ _06753_ VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__xor2_2
X_18914_ _11310_ _11312_ VGND VGND VPWR VPWR _11337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19894_ _01691_ _01708_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18845_ _11263_ _11269_ VGND VGND VPWR VPWR _11270_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_235_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18776_ _11191_ _11185_ _11202_ VGND VGND VPWR VPWR _11204_ sky130_fd_sc_hd__nand3_1
XTAP_5690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15988_ _08152_ _08353_ _08558_ VGND VGND VPWR VPWR _08597_ sky130_fd_sc_hd__o21a_1
XFILLER_0_222_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17727_ _10234_ _10235_ VGND VGND VPWR VPWR _10236_ sky130_fd_sc_hd__nor2_4
XFILLER_0_89_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14939_ _07608_ _05735_ _07609_ _07092_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__o211a_1
Xclkbuf_4_11__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_4_11__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17658_ top_inst.grid_inst.data_path_wires\[11\]\[1\] top_inst.grid_inst.data_path_wires\[11\]\[0\]
+ _10056_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _10169_ sky130_fd_sc_hd__and4_1
XFILLER_0_77_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16609_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[16\] _07866_ VGND
+ VGND VPWR VPWR _09183_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17589_ _10100_ _10101_ _10085_ VGND VGND VPWR VPWR _10103_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_15_clk clknet_4_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19328_ _04873_ VGND VGND VPWR VPWR _11722_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19259_ _11635_ _11658_ VGND VGND VPWR VPWR _11673_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_1291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22270_ _03709_ _03686_ _03906_ _03957_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21221_ _07707_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__buf_4
Xhold100 top_inst.deskew_buff_inst.col_input\[66\] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold111 _00283_ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold122 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[29\] VGND
+ VGND VPWR VPWR net304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold133 top_inst.deskew_buff_inst.col_input\[46\] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold144 _00040_ VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__dlygate4sd3_1
X_21152_ _02897_ _02021_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__or2_1
Xhold155 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[7\] VGND
+ VGND VPWR VPWR net337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold166 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[4\] VGND
+ VGND VPWR VPWR net348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold177 top_inst.axis_out_inst.out_buff_data\[14\] VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20103_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[27\] _01761_ _01762_
+ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__a21o_1
Xhold188 _00290_ VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _00940_ VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21083_ _02832_ _02833_ _02830_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20034_ _01845_ _01849_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__xor2_2
XFILLER_0_77_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21985_ _02873_ _02877_ _03692_ _03660_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__o211a_1
XFILLER_0_241_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23724_ clknet_leaf_120_clk _00257_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20936_ _04868_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__buf_6
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23655_ clknet_leaf_135_clk _00188_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_20867_ _01819_ _02637_ _02639_ _02035_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22606_ _04248_ _04251_ _04277_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_119_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_942 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23586_ clknet_leaf_106_clk net271 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_20798_ _02462_ _02554_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22537_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[16\] _04215_ _04216_
+ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13270_ _06044_ _06045_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22468_ _04149_ _04150_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__and2_1
XFILLER_0_224_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24207_ clknet_leaf_17_clk _00740_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_12221_ _05127_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__buf_2
X_21419_ _03118_ _03119_ _03153_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__and3_1
X_22399_ _04055_ _04056_ _04082_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__nand3_1
XFILLER_0_20_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12152_ net741 _05097_ _05100_ _05101_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__o211a_1
X_24138_ clknet_leaf_144_clk _00671_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_1004 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16960_ _09470_ _09472_ _09471_ VGND VGND VPWR VPWR _09515_ sky130_fd_sc_hd__a21bo_1
X_12083_ net546 _05058_ _05061_ _05062_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24069_ clknet_leaf_84_clk _00602_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15911_ _08517_ _08521_ VGND VGND VPWR VPWR _08522_ sky130_fd_sc_hd__xor2_1
XFILLER_0_235_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16891_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[7\] _09397_ _09396_
+ VGND VGND VPWR VPWR _09448_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18630_ _11042_ _11064_ _11062_ VGND VGND VPWR VPWR _11089_ sky130_fd_sc_hd__o21a_1
XFILLER_0_216_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15842_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[10\] _08374_ VGND
+ VGND VPWR VPWR _08455_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_217_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18561_ _10933_ _11020_ VGND VGND VPWR VPWR _11022_ sky130_fd_sc_hd__or2_1
XFILLER_0_232_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _08335_ _08337_ VGND VGND VPWR VPWR _08388_ sky130_fd_sc_hd__and2b_1
XFILLER_0_235_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12985_ _05772_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__clkbuf_4
XTAP_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17512_ _10030_ _09215_ VGND VGND VPWR VPWR _10039_ sky130_fd_sc_hd__or2_2
XTAP_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14724_ _07079_ _07074_ _07089_ VGND VGND VPWR VPWR _07412_ sky130_fd_sc_hd__and3_1
XTAP_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ top_inst.axis_out_inst.out_buff_data\[41\] _04969_ VGND VGND VPWR VPWR _04978_
+ sky130_fd_sc_hd__or2_1
X_18492_ _10911_ _10954_ VGND VGND VPWR VPWR _10955_ sky130_fd_sc_hd__xnor2_1
XTAP_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17443_ _09978_ _09979_ VGND VGND VPWR VPWR _09980_ sky130_fd_sc_hd__or2_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14655_ _07342_ _07343_ _07325_ VGND VGND VPWR VPWR _07345_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[11\] _04930_
+ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__or2_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1028 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13606_ _06273_ _06311_ _06309_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__a21o_1
X_17374_ _09624_ _09912_ VGND VGND VPWR VPWR _09914_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14586_ _07070_ _07082_ _07239_ _07238_ VGND VGND VPWR VPWR _07277_ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11798_ net856 _04898_ _04899_ _04889_ VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19113_ _11482_ _11484_ _11486_ VGND VGND VPWR VPWR _11532_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16325_ _08845_ _08854_ _08906_ VGND VGND VPWR VPWR _08907_ sky130_fd_sc_hd__o21a_1
XFILLER_0_137_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13537_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[5\] _06242_ _06285_
+ _06286_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19044_ _11463_ _11464_ VGND VGND VPWR VPWR _11465_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16256_ top_inst.grid_inst.data_path_wires\[8\]\[4\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[3\]
+ top_inst.grid_inst.data_path_wires\[8\]\[3\] _08693_ VGND VGND VPWR VPWR _08839_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13468_ _05317_ _06221_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__nand2_1
XFILLER_0_207_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15207_ _07793_ _07802_ _07854_ VGND VGND VPWR VPWR _07855_ sky130_fd_sc_hd__o21a_1
X_12419_ net286 _05243_ _05253_ _05247_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__o211a_1
X_16187_ _08750_ _08753_ _08751_ VGND VGND VPWR VPWR _08772_ sky130_fd_sc_hd__o21ai_1
X_13399_ _06161_ _06164_ _06098_ VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15138_ top_inst.grid_inst.data_path_wires\[6\]\[3\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[6\]\[4\]
+ VGND VGND VPWR VPWR _07787_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19946_ _01561_ _01765_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__nor2_1
X_15069_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[4\] _07689_ _07690_
+ VGND VGND VPWR VPWR _07720_ sky130_fd_sc_hd__a21boi_2
Xclkbuf_leaf_4_clk clknet_4_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19877_ _01528_ _01699_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__xor2_2
XFILLER_0_177_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18828_ _11229_ _11253_ VGND VGND VPWR VPWR _11254_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18759_ _11175_ _11187_ VGND VGND VPWR VPWR _11188_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21770_ _03246_ _03492_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__and2_1
XFILLER_0_176_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20721_ _02496_ _02497_ _02466_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_1076 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23440_ top_inst.axis_out_inst.out_buff_data\[108\] _04835_ VGND VGND VPWR VPWR _04842_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_50_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20652_ _02430_ _02431_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23371_ _04684_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20583_ _02241_ _02328_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__or2b_2
XFILLER_0_2_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22322_ _04005_ _04007_ _05311_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22253_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[9\] _03894_ VGND
+ VGND VPWR VPWR _03941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21204_ _02871_ _02868_ _02885_ _02882_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__nand4_1
XFILLER_0_197_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22184_ _03859_ _03873_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21135_ _02864_ _02881_ _02886_ _02880_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21066_ _02503_ _02812_ _02793_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_217_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20017_ _01809_ _01826_ _01833_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__a21o_1
XFILLER_0_214_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_1220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12770_ _05564_ _05540_ _05578_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21968_ _03680_ _02869_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23707_ clknet_leaf_124_clk _00240_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20919_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[23\] _02467_ VGND
+ VGND VPWR VPWR _02689_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21899_ _03596_ _03616_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_167_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _07135_ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__clkbuf_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23638_ clknet_leaf_108_clk net399 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14371_ _05772_ VGND VGND VPWR VPWR _07075_ sky130_fd_sc_hd__buf_2
XFILLER_0_135_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23569_ clknet_leaf_103_clk _00102_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16110_ _08683_ _08661_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _08700_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13322_ _06016_ net182 _06096_ VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_51_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17090_ _09553_ _09640_ _09641_ VGND VGND VPWR VPWR _09642_ sky130_fd_sc_hd__or3_1
XFILLER_0_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_243_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16041_ _08626_ _08648_ _04870_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__o21a_1
X_13253_ _05986_ _05991_ _06029_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_1224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12204_ net895 _05123_ _05131_ _05128_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__o211a_1
X_13184_ _05925_ _05921_ _05962_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_1292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19800_ _01596_ _01620_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__nor2_1
X_12135_ net820 _05089_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__or2_1
X_17992_ _10490_ _10494_ VGND VGND VPWR VPWR _10495_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16943_ _09462_ _09461_ VGND VGND VPWR VPWR _09498_ sky130_fd_sc_hd__and2b_1
X_19731_ _01518_ _01556_ _01554_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12066_ net717 _05050_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__or2_1
XFILLER_0_236_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16874_ _09428_ _09429_ _09430_ VGND VGND VPWR VPWR _09431_ sky130_fd_sc_hd__nand3_1
X_19662_ _01489_ _01490_ _01491_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__nand3_1
XFILLER_0_204_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15825_ _08163_ _08169_ _08353_ _08143_ VGND VGND VPWR VPWR _08438_ sky130_fd_sc_hd__o2bb2a_1
X_18613_ _10071_ _11071_ _11072_ _10620_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_205_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19593_ _01422_ _01423_ _01392_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__a21o_1
XTAP_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15756_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[1\] _08154_ top_inst.grid_inst.data_path_wires\[7\]\[7\]
+ VGND VGND VPWR VPWR _08371_ sky130_fd_sc_hd__o21ai_2
X_18544_ _10967_ _10973_ _10971_ VGND VGND VPWR VPWR _11005_ sky130_fd_sc_hd__a21o_1
XTAP_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12968_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _05761_ sky130_fd_sc_hd__clkbuf_4
XTAP_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14707_ _07361_ _07362_ _07394_ _07395_ VGND VGND VPWR VPWR _07396_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_87_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11919_ net1001 _04964_ _04967_ _04968_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18475_ _10592_ _10610_ _10934_ _10937_ VGND VGND VPWR VPWR _10938_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15687_ _08302_ _08303_ VGND VGND VPWR VPWR _08304_ sky130_fd_sc_hd__nor2_1
XFILLER_0_213_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12899_ _05701_ _05703_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__nor2_1
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _09919_ _09918_ _09937_ _09940_ VGND VGND VPWR VPWR _09964_ sky130_fd_sc_hd__o31a_1
XFILLER_0_185_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14638_ _07070_ _07090_ VGND VGND VPWR VPWR _07328_ sky130_fd_sc_hd__nand2_4
XFILLER_0_184_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17357_ _09896_ _09897_ VGND VGND VPWR VPWR _09898_ sky130_fd_sc_hd__and2b_1
X_14569_ _07258_ _07259_ _07260_ VGND VGND VPWR VPWR _07261_ sky130_fd_sc_hd__or3_4
XFILLER_0_166_1015 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16308_ _08838_ _08841_ _08842_ VGND VGND VPWR VPWR _08890_ sky130_fd_sc_hd__and3_1
XFILLER_0_141_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17288_ _09625_ _09814_ VGND VGND VPWR VPWR _09832_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19027_ _11446_ _11447_ VGND VGND VPWR VPWR _11448_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16239_ _08820_ _08821_ _08792_ _08793_ VGND VGND VPWR VPWR _08823_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_28_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_535 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19929_ _01709_ _01732_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_215_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22940_ net404 _04557_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__or2_1
XFILLER_0_177_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22871_ net762 _04509_ _04518_ _04511_ VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24610_ clknet_leaf_21_clk _01143_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_218_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21822_ _03510_ _03523_ _03542_ _01984_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__a31o_1
XFILLER_0_223_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24541_ clknet_leaf_102_clk _01074_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21753_ _03473_ _03477_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20704_ _02459_ _02482_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__xnor2_1
X_24472_ clknet_leaf_55_clk _01005_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_1172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21684_ _03403_ _03411_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23423_ net371 _04827_ _04832_ _04831_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20635_ _02391_ _02392_ _02415_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23354_ net473 _04791_ _04794_ _04795_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20566_ _02135_ _02348_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22305_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[18\]\[3\]
+ _03953_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__and3_1
XFILLER_0_171_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23285_ net489 _04752_ _04755_ _04756_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__o211a_1
X_20497_ _02275_ _02280_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22236_ _03713_ _03878_ _03924_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_225_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22167_ _03850_ _03856_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21118_ _02873_ _02869_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_1016 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22098_ _03788_ _03789_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__nand2_1
XFILLER_0_218_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1038 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13940_ _06624_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[1\] _06622_
+ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _06661_ sky130_fd_sc_hd__nand4_2
X_21049_ _02812_ _02813_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__or2_1
XFILLER_0_227_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13871_ _06496_ _06591_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__nor2_1
XFILLER_0_242_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15610_ _08226_ _08228_ VGND VGND VPWR VPWR _08229_ sky130_fd_sc_hd__xor2_2
XFILLER_0_236_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12822_ _05591_ _05593_ _05628_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__or3_1
X_16590_ _09137_ _09139_ _09163_ _09164_ VGND VGND VPWR VPWR _09165_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_9_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_243_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_232_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15541_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _08167_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12753_ _05552_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18260_ top_inst.grid_inst.data_path_wires\[12\]\[2\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[12\]\[3\]
+ VGND VGND VPWR VPWR _10728_ sky130_fd_sc_hd__a22oi_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15472_ _08086_ _08087_ _08084_ VGND VGND VPWR VPWR _08113_ sky130_fd_sc_hd__o21a_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12684_ _05448_ _05452_ _05450_ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_38_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _09735_ _09758_ VGND VGND VPWR VPWR _09759_ sky130_fd_sc_hd__xnor2_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14423_ _07066_ _07069_ _07073_ _07062_ VGND VGND VPWR VPWR _07119_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18191_ _05887_ _10659_ _10660_ _10661_ VGND VGND VPWR VPWR _10662_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17142_ _06140_ _09692_ VGND VGND VPWR VPWR _09693_ sky130_fd_sc_hd__nand2_1
X_14354_ _07060_ VGND VGND VPWR VPWR _07061_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13305_ _06073_ _06075_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17073_ _09624_ VGND VGND VPWR VPWR _09625_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_150_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14285_ _06978_ VGND VGND VPWR VPWR _06995_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16024_ _08629_ _08631_ VGND VGND VPWR VPWR _08632_ sky130_fd_sc_hd__xnor2_1
X_13236_ _06011_ _06012_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13167_ _05904_ _05945_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12118_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[23\] _05076_
+ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13098_ _05874_ _05875_ _05878_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__nor3_1
XFILLER_0_104_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17975_ _10477_ _10478_ VGND VGND VPWR VPWR _10479_ sky130_fd_sc_hd__or2_1
XFILLER_0_236_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19714_ _01488_ _01496_ _01495_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_40_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16926_ _09478_ _09479_ _09480_ VGND VGND VPWR VPWR _09482_ sky130_fd_sc_hd__a21o_1
X_12049_ net919 _05031_ _05042_ _05035_ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19645_ _01438_ _01437_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__and2b_1
X_16857_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[7\] _09364_ _09365_
+ VGND VGND VPWR VPWR _09414_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_204_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15808_ _08368_ _08366_ VGND VGND VPWR VPWR _08422_ sky130_fd_sc_hd__and2b_1
X_16788_ _09344_ _09345_ _09311_ VGND VGND VPWR VPWR _09347_ sky130_fd_sc_hd__a21oi_1
X_19576_ _01297_ _01314_ _11686_ net239 VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__or4b_4
XFILLER_0_88_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15739_ top_inst.grid_inst.data_path_wires\[7\]\[2\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[6\]
+ _08353_ top_inst.grid_inst.data_path_wires\[7\]\[1\] VGND VGND VPWR VPWR _08354_
+ sky130_fd_sc_hd__o2bb2a_1
X_18527_ _10986_ _10988_ VGND VGND VPWR VPWR _10989_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18458_ _10887_ _10886_ VGND VGND VPWR VPWR _10921_ sky130_fd_sc_hd__or2b_1
XFILLER_0_29_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17409_ _05405_ _09947_ VGND VGND VPWR VPWR _09948_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18389_ _10852_ _10853_ VGND VGND VPWR VPWR _10854_ sky130_fd_sc_hd__xor2_1
XFILLER_0_117_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20420_ _02160_ _02162_ _02204_ _02205_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_172_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_244_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20351_ _01992_ _02015_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[6\]
+ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23070_ top_inst.axis_in_inst.inbuf_bus\[22\] _04629_ VGND VGND VPWR VPWR _04633_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_114_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20282_ top_inst.deskew_buff_inst.col_input\[35\] _05730_ VGND VGND VPWR VPWR _02072_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_222_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22021_ net1014 _06169_ _03717_ _03702_ VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23972_ clknet_leaf_114_clk _00505_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22923_ net1029 _04535_ _04547_ _04537_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_233_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22854_ net1039 _04496_ _04508_ _04498_ VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21805_ _03527_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22785_ _04452_ _04453_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24524_ clknet_leaf_131_clk _01057_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dfxtp_2
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21736_ _03460_ _03461_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__nor2_2
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24455_ clknet_leaf_54_clk _00988_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_21667_ _03340_ _03395_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23406_ net751 _04655_ _04823_ _04819_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20618_ _02397_ _02398_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__nand2_1
X_24386_ clknet_leaf_38_clk _00919_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_978 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21598_ _03325_ _03326_ _03328_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_151_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23337_ top_inst.axis_out_inst.out_buff_data\[94\] _04778_ _04785_ _04782_ VGND VGND
+ VPWR VPWR _01118_ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20549_ _02331_ _02288_ _02289_ _02241_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14070_ top_inst.grid_inst.data_path_wires\[3\]\[6\] _06785_ VGND VGND VPWR VPWR
+ _06786_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23268_ net776 _04739_ _04746_ _04743_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13021_ top_inst.grid_inst.data_path_wires\[1\]\[4\] top_inst.grid_inst.data_path_wires\[1\]\[3\]
+ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__nand4_1
XFILLER_0_131_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22219_ _03711_ top_inst.grid_inst.data_path_wires\[18\]\[1\] _03868_ VGND VGND VPWR
+ VPWR _03908_ sky130_fd_sc_hd__and3_1
XFILLER_0_219_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23199_ net789 _04700_ _04707_ _04704_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__o211a_1
XTAP_6721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14972_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _07633_ sky130_fd_sc_hd__clkbuf_4
X_17760_ _10266_ _10268_ VGND VGND VPWR VPWR _10269_ sky130_fd_sc_hd__nor2_1
XFILLER_0_233_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16711_ _09270_ _09271_ VGND VGND VPWR VPWR _09272_ sky130_fd_sc_hd__and2_1
X_13923_ _06628_ _06647_ _06649_ _06639_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17691_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[7\] _10200_ VGND
+ VGND VPWR VPWR _10201_ sky130_fd_sc_hd__xor2_2
XFILLER_0_215_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16642_ _09209_ VGND VGND VPWR VPWR _09210_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19430_ net231 _01263_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[6\]
+ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_187_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13854_ _06593_ _06594_ VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__nor2_1
XFILLER_0_202_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12805_ _05571_ _05572_ _05612_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16573_ _09148_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__clkbuf_1
X_19361_ top_inst.deskew_buff_inst.col_input\[3\] _05730_ VGND VGND VPWR VPWR _01199_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_29_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13785_ _06525_ _06526_ _06527_ VGND VGND VPWR VPWR _06528_ sky130_fd_sc_hd__o21a_1
XFILLER_0_186_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15524_ _08154_ VGND VGND VPWR VPWR _08155_ sky130_fd_sc_hd__clkbuf_4
X_18312_ _10777_ _10778_ VGND VGND VPWR VPWR _10779_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_210_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12736_ _05497_ _05500_ _05498_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__o21ba_1
X_19292_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _11693_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_155_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _10683_ _10699_ VGND VGND VPWR VPWR _10711_ sky130_fd_sc_hd__nand2_1
XFILLER_0_210_1266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15455_ _08094_ _08095_ _05315_ VGND VGND VPWR VPWR _08097_ sky130_fd_sc_hd__o21a_1
X_12667_ _05435_ _05437_ _05476_ _05477_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_26_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14406_ _07066_ _07065_ _07069_ _07062_ VGND VGND VPWR VPWR _07103_ sky130_fd_sc_hd__a22o_1
XFILLER_0_203_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18174_ top_inst.grid_inst.data_path_wires\[12\]\[1\] top_inst.grid_inst.data_path_wires\[12\]\[0\]
+ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _10645_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15386_ net974 _05403_ VGND VGND VPWR VPWR _08029_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12598_ _05383_ _05410_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17125_ _09674_ _09675_ _09551_ _09552_ VGND VGND VPWR VPWR _09676_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14337_ _07043_ _07044_ _05633_ VGND VGND VPWR VPWR _07046_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold507 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[30\] VGND
+ VGND VPWR VPWR net689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold518 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[23\] VGND
+ VGND VPWR VPWR net700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17056_ _09594_ _09607_ _09608_ VGND VGND VPWR VPWR _09609_ sky130_fd_sc_hd__and3_1
Xhold529 top_inst.deskew_buff_inst.col_input\[107\] VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14268_ _06977_ _06898_ _06934_ VGND VGND VPWR VPWR _06979_ sky130_fd_sc_hd__or3_2
XFILLER_0_180_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_1436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16007_ _08578_ _08579_ _08615_ VGND VGND VPWR VPWR _08616_ sky130_fd_sc_hd__a21boi_2
X_13219_ _05950_ _05996_ _05947_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14199_ _06866_ _06871_ _06911_ VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__a21oi_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1002 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _10460_ _10461_ VGND VGND VPWR VPWR _10462_ sky130_fd_sc_hd__and2_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16909_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[2\] _09218_ VGND
+ VGND VPWR VPWR _09465_ sky130_fd_sc_hd__nand2_2
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17889_ _10352_ _10327_ VGND VGND VPWR VPWR _10395_ sky130_fd_sc_hd__or2b_1
XFILLER_0_205_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19628_ _01456_ _01457_ _01440_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_672 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19559_ _01355_ _01351_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__and2b_1
XFILLER_0_215_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22570_ _04225_ _04247_ _04238_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21521_ top_inst.grid_inst.data_path_wires\[17\]\[5\] _02897_ VGND VGND VPWR VPWR
+ _03254_ sky130_fd_sc_hd__and2b_1
XFILLER_0_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24240_ clknet_leaf_113_clk _00773_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_113_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21452_ _03184_ _03186_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__xor2_2
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20403_ _02186_ _02187_ _02188_ _01989_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__a22o_1
X_24171_ clknet_leaf_23_clk _00704_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21383_ _03104_ _03074_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__or2b_1
XFILLER_0_86_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23122_ net88 _04659_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__or2_1
XFILLER_0_226_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20334_ _02104_ _02105_ _02120_ _02121_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23053_ net971 _04616_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__or2_1
Xoutput38 net38 VGND VGND VPWR VPWR output_tdata[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20265_ _01992_ _02009_ _02052_ _02053_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput49 net49 VGND VGND VPWR VPWR output_tdata[10] sky130_fd_sc_hd__clkbuf_4
XTAP_6017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22004_ _03705_ _05275_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__or2_1
XTAP_6039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20196_ _04858_ _11700_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__or2_2
XTAP_5316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_215_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23955_ clknet_leaf_91_clk _00488_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22906_ net396 _04535_ _04538_ _04537_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23886_ clknet_leaf_64_clk _00419_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_233_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22837_ net655 _04496_ _04499_ _04498_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13570_ _06263_ _06317_ _06318_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__a21oi_1
X_22768_ _04436_ _04437_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ net1005 _05314_ _05337_ _05308_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24507_ clknet_leaf_132_clk _01040_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dfxtp_2
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21719_ _03441_ _03438_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__or2b_1
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22699_ _04092_ _04370_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__nand2_1
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15240_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[8\] _07845_ _07844_
+ VGND VGND VPWR VPWR _07887_ sky130_fd_sc_hd__a21o_1
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24438_ clknet_leaf_57_clk _00971_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12452_ top_inst.skew_buff_inst.row\[0\].output_reg\[1\] top_inst.axis_in_inst.inbuf_bus\[1\]
+ net211 VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__mux2_2
XFILLER_0_124_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15171_ _07771_ _07811_ VGND VGND VPWR VPWR _07819_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24369_ clknet_leaf_37_clk net937 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].output_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12383_ net373 _05222_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14122_ _06789_ _06783_ VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__or2b_1
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14053_ _06742_ _06747_ VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__nor2_1
X_18930_ _11350_ _11352_ VGND VGND VPWR VPWR _11353_ sky130_fd_sc_hd__and2b_1
XFILLER_0_240_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13004_ _05787_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__buf_4
XFILLER_0_219_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18861_ _11260_ _11261_ _11284_ _11285_ VGND VGND VPWR VPWR _11286_ sky130_fd_sc_hd__a211oi_2
XTAP_6540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17812_ _10279_ _10319_ VGND VGND VPWR VPWR _10320_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_219_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18792_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[13\]\[1\]
+ top_inst.grid_inst.data_path_wires\[13\]\[0\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[4\]
+ VGND VGND VPWR VPWR _11219_ sky130_fd_sc_hd__a22o_1
XTAP_6595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14955_ top_inst.grid_inst.data_path_wires\[6\]\[6\] VGND VGND VPWR VPWR _07621_
+ sky130_fd_sc_hd__buf_2
X_17743_ _10027_ _10054_ _10213_ _10251_ VGND VGND VPWR VPWR _10252_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_89_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13906_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _06637_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14886_ _07540_ _07544_ _07569_ VGND VGND VPWR VPWR _07570_ sky130_fd_sc_hd__a21o_1
X_17674_ _10182_ _10183_ _10154_ _10155_ VGND VGND VPWR VPWR _10185_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_187_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19413_ _01207_ _01210_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__nand2_1
X_16625_ top_inst.skew_buff_inst.row\[2\].output_reg\[2\] top_inst.axis_in_inst.inbuf_bus\[18\]
+ _07059_ VGND VGND VPWR VPWR _09196_ sky130_fd_sc_hd__mux2_4
XFILLER_0_202_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13837_ _06575_ _06577_ VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_806 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_202_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16556_ _09125_ _09131_ VGND VGND VPWR VPWR _09132_ sky130_fd_sc_hd__xnor2_1
X_19344_ _11729_ _11730_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__or2_1
X_13768_ _06510_ _06511_ VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12719_ _05447_ _05449_ _05283_ _05528_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__or4_1
X_15507_ top_inst.grid_inst.data_path_wires\[7\]\[3\] VGND VGND VPWR VPWR _08143_
+ sky130_fd_sc_hd__buf_4
X_16487_ _09021_ _09024_ _09064_ VGND VGND VPWR VPWR _09065_ sky130_fd_sc_hd__a21bo_1
X_19275_ _11678_ VGND VGND VPWR VPWR _11679_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_155_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_13699_ _06443_ _06444_ _05328_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15438_ _08005_ _08078_ VGND VGND VPWR VPWR _08080_ sky130_fd_sc_hd__and2_1
X_18226_ _10693_ _10694_ VGND VGND VPWR VPWR _10695_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_870 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15369_ _08011_ _08012_ VGND VGND VPWR VPWR _08013_ sky130_fd_sc_hd__xnor2_1
X_18157_ _10599_ _10600_ _10597_ _10581_ VGND VGND VPWR VPWR _10629_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17108_ _09621_ _09658_ _09292_ VGND VGND VPWR VPWR _09660_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold304 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[18\] VGND
+ VGND VPWR VPWR net486 sky130_fd_sc_hd__dlygate4sd3_1
X_18088_ _10577_ _08674_ VGND VGND VPWR VPWR _10578_ sky130_fd_sc_hd__or2_1
Xhold315 top_inst.deskew_buff_inst.col_input\[36\] VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 top_inst.deskew_buff_inst.col_input\[112\] VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold337 _00134_ VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold348 top_inst.axis_out_inst.out_buff_data\[127\] VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__dlygate4sd3_1
X_17039_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[12\] _09419_ VGND
+ VGND VPWR VPWR _09592_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold359 top_inst.axis_out_inst.out_buff_data\[6\] VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20050_ _01837_ _01860_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23740_ clknet_leaf_127_clk _00273_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20952_ _02718_ _02719_ _02473_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_178_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23671_ clknet_leaf_116_clk net813 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_20883_ _02653_ _02654_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22622_ _04275_ _04298_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22553_ _04231_ _04232_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21504_ _03198_ _03197_ _03230_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_174_894 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22484_ _04061_ _04165_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24223_ clknet_leaf_19_clk _00756_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21435_ _02875_ _03168_ _03169_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_146_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24154_ clknet_leaf_18_clk _00687_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21366_ _03043_ _03057_ _03102_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__o21a_1
XFILLER_0_142_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23105_ net331 _05323_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__or2_1
X_20317_ _02102_ _02103_ _02089_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__a21oi_1
X_24085_ clknet_leaf_87_clk _00618_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold860 top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[15\] VGND VGND
+ VPWR VPWR net1042 sky130_fd_sc_hd__dlygate4sd3_1
X_21297_ _03007_ _03016_ _03018_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__o21ai_1
Xhold871 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[4\] VGND VGND
+ VPWR VPWR net1053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[1\] VGND VGND
+ VPWR VPWR net1064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23036_ net606 _04603_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__or2_1
Xhold893 top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[0\] VGND VGND
+ VPWR VPWR net1075 sky130_fd_sc_hd__dlygate4sd3_1
X_20248_ _01993_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[0\] VGND
+ VGND VPWR VPWR _02039_ sky130_fd_sc_hd__and2_1
XTAP_5102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20179_ _10030_ _11677_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__or2_1
XTAP_5146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_216_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14740_ _07409_ _07427_ VGND VGND VPWR VPWR _07428_ sky130_fd_sc_hd__or2_1
XTAP_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23938_ clknet_leaf_81_clk _00471_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ net553 _04982_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14671_ _07350_ _07353_ VGND VGND VPWR VPWR _07360_ sky130_fd_sc_hd__nand2_1
XTAP_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23869_ clknet_leaf_78_clk _00402_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[18\] _04943_
+ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__or2_1
XFILLER_0_233_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16410_ _08952_ _08989_ VGND VGND VPWR VPWR _08990_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13622_ _06367_ _06368_ VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__nor2_1
X_17390_ _09905_ _09926_ VGND VGND VPWR VPWR _09929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16341_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[8\]\[3\]
+ top_inst.grid_inst.data_path_wires\[8\]\[2\] _08876_ VGND VGND VPWR VPWR _08922_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_27_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13553_ _06300_ _06301_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12504_ _05318_ _05321_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19060_ _11140_ _11143_ _11164_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _11480_ sky130_fd_sc_hd__and4b_1
X_16272_ _08845_ _08854_ VGND VGND VPWR VPWR _08855_ sky130_fd_sc_hd__xor2_1
X_13484_ _06233_ _06234_ _06235_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__and3b_1
XFILLER_0_124_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15223_ top_inst.grid_inst.data_path_wires\[6\]\[2\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[7\]
+ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[6\]\[3\]
+ VGND VGND VPWR VPWR _07870_ sky130_fd_sc_hd__and4b_1
XFILLER_0_125_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18011_ _10473_ _10512_ _10513_ VGND VGND VPWR VPWR _10514_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12435_ net335 _05256_ _05263_ _05261_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15154_ _07793_ _07802_ VGND VGND VPWR VPWR _07803_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12366_ net432 _05222_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__or2_1
XFILLER_0_239_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14105_ _06814_ _06819_ VGND VGND VPWR VPWR _06820_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19962_ _01561_ _01780_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__xor2_2
X_15085_ _07709_ _07735_ VGND VGND VPWR VPWR _07736_ sky130_fd_sc_hd__nand2_1
X_12297_ net456 _05183_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__or2_1
X_14036_ _06751_ _06752_ VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__nor2_1
X_18913_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[7\] _11302_ _11303_
+ VGND VGND VPWR VPWR _11336_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_120_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19893_ _01691_ _01708_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18844_ _11264_ _11268_ VGND VGND VPWR VPWR _11269_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18775_ _11191_ _11185_ _11202_ VGND VGND VPWR VPWR _11203_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15987_ _08517_ _08559_ _08560_ VGND VGND VPWR VPWR _08596_ sky130_fd_sc_hd__o21ba_1
XTAP_5691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17726_ top_inst.grid_inst.data_path_wires\[11\]\[7\] _10044_ _10042_ VGND VGND VPWR
+ VPWR _10235_ sky130_fd_sc_hd__and3_1
XFILLER_0_188_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14938_ _05739_ _07292_ VGND VGND VPWR VPWR _07609_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17657_ _10022_ _10056_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[5\]
+ _10025_ VGND VGND VPWR VPWR _10168_ sky130_fd_sc_hd__a22oi_1
X_14869_ _07550_ _07552_ VGND VGND VPWR VPWR _07554_ sky130_fd_sc_hd__or2_1
XFILLER_0_159_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_230_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16608_ _09165_ _09167_ _09168_ _09181_ VGND VGND VPWR VPWR _09182_ sky130_fd_sc_hd__o31a_1
XFILLER_0_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17588_ _10085_ _10100_ _10101_ VGND VGND VPWR VPWR _10102_ sky130_fd_sc_hd__or3_1
XFILLER_0_175_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19327_ net932 _10616_ _11721_ _11714_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__o211a_1
X_16539_ _09079_ _09115_ _04867_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19258_ _11663_ _11671_ VGND VGND VPWR VPWR _11672_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18209_ _10656_ _10659_ VGND VGND VPWR VPWR _10679_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_1224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19189_ _11596_ _11605_ VGND VGND VPWR VPWR _11606_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21220_ _02958_ _02959_ _07595_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__a21o_1
Xhold101 _00041_ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[6\] VGND VGND
+ VPWR VPWR net294 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold123 _00292_ VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 _00117_ VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold145 top_inst.deskew_buff_inst.col_input\[61\] VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__buf_1
X_21151_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _02897_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_229_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold156 _00014_ VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 _00011_ VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20102_ _01891_ _01894_ _01893_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__a21o_1
Xhold178 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[6\] VGND
+ VGND VPWR VPWR net360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 top_inst.deskew_buff_inst.col_input\[100\] VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__dlygate4sd3_1
X_21082_ _02844_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20033_ _01847_ _01848_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21984_ _03690_ _03691_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__or2_1
XFILLER_0_240_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23723_ clknet_leaf_120_clk _00256_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20935_ net647 _02638_ VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__or2_1
XFILLER_0_230_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23654_ clknet_leaf_135_clk _00187_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20866_ net861 _02638_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22605_ _04253_ _04255_ _04278_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__nand3_1
XFILLER_0_7_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23585_ clknet_leaf_106_clk net279 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20797_ _02558_ _02560_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__nand2_1
XFILLER_0_221_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22536_ _03938_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22467_ _04124_ _04125_ _04148_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__nand3_1
XFILLER_0_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12220_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[3\] _05129_
+ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__or2_1
X_24206_ clknet_leaf_117_clk _00739_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_21418_ _03118_ _03119_ _03153_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_103_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22398_ _04055_ _04056_ _04082_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12151_ _04994_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__clkbuf_4
X_24137_ clknet_leaf_144_clk _00670_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21349_ _03084_ _03085_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24068_ clknet_leaf_84_clk _00601_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_12082_ _04994_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__buf_2
Xhold690 top_inst.axis_out_inst.out_buff_data\[103\] VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1016 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23019_ net903 _04603_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15910_ _08519_ _08520_ VGND VGND VPWR VPWR _08521_ sky130_fd_sc_hd__or2_1
X_16890_ _09410_ net183 VGND VGND VPWR VPWR _09447_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _08152_ _08159_ _08405_ _08406_ VGND VGND VPWR VPWR _08454_ sky130_fd_sc_hd__a31o_1
XFILLER_0_244_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_232_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ _10933_ _11020_ VGND VGND VPWR VPWR _11021_ sky130_fd_sc_hd__nand2_1
XTAP_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _05274_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__buf_4
XTAP_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ _08385_ _08386_ VGND VGND VPWR VPWR _08387_ sky130_fd_sc_hd__xnor2_1
XTAP_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17511_ _10037_ VGND VGND VPWR VPWR _10038_ sky130_fd_sc_hd__clkbuf_4
XTAP_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14723_ _07377_ _07385_ VGND VGND VPWR VPWR _07411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11935_ _04911_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__clkbuf_4
XTAP_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18491_ _10952_ _10953_ VGND VGND VPWR VPWR _10954_ sky130_fd_sc_hd__and2_1
XTAP_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14654_ _07325_ _07342_ _07343_ VGND VGND VPWR VPWR _07344_ sky130_fd_sc_hd__nand3_1
X_17442_ _09977_ _09972_ VGND VGND VPWR VPWR _09979_ sky130_fd_sc_hd__and2b_1
XFILLER_0_68_951 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _04911_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__clkbuf_4
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13605_ _06350_ _06352_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14585_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[7\] _07230_ _07229_
+ _07066_ VGND VGND VPWR VPWR _07276_ sky130_fd_sc_hd__a22o_1
X_17373_ _09624_ _09912_ VGND VGND VPWR VPWR _09913_ sky130_fd_sc_hd__or2_2
XFILLER_0_32_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11797_ net468 _04890_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19112_ _11529_ _11530_ VGND VGND VPWR VPWR _11531_ sky130_fd_sc_hd__nand2_1
X_16324_ _08832_ _08844_ VGND VGND VPWR VPWR _08906_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13536_ _06259_ _06284_ _05399_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16255_ _08798_ _08837_ VGND VGND VPWR VPWR _08838_ sky130_fd_sc_hd__xor2_1
X_19043_ _11427_ _11462_ VGND VGND VPWR VPWR _11464_ sky130_fd_sc_hd__or2_1
X_13467_ _06217_ _06219_ _06220_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15206_ _07780_ _07792_ VGND VGND VPWR VPWR _07854_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12418_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[24\] _05248_
+ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__or2_1
XFILLER_0_242_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16186_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[4\] _08743_ _08744_
+ VGND VGND VPWR VPWR _08771_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13398_ _06098_ _06161_ _06164_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15137_ _07746_ _07785_ VGND VGND VPWR VPWR _07786_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12349_ net288 _05209_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19945_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[21\] _01764_ VGND
+ VGND VPWR VPWR _01765_ sky130_fd_sc_hd__xnor2_1
X_15068_ _07717_ _07718_ VGND VGND VPWR VPWR _07719_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14019_ _06715_ _06720_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19876_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[18\] _01480_ VGND
+ VGND VPWR VPWR _01699_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_208_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18827_ _11250_ _11252_ VGND VGND VPWR VPWR _11253_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_235_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18758_ _11185_ _11186_ VGND VGND VPWR VPWR _11187_ sky130_fd_sc_hd__and2_1
XFILLER_0_222_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17709_ _10195_ _10218_ VGND VGND VPWR VPWR _10219_ sky130_fd_sc_hd__xor2_1
XFILLER_0_222_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18689_ _10599_ _10584_ _11134_ _10620_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20720_ _02466_ _02496_ _02497_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__and3_1
XFILLER_0_172_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20651_ _02004_ _02016_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[13\]
+ VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23370_ net714 _04791_ _04803_ _04795_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20582_ _02009_ _02329_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__and2_2
XFILLER_0_74_998 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22321_ _04005_ _04007_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22252_ _03898_ _03901_ _03899_ VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_60_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21203_ top_inst.grid_inst.data_path_wires\[17\]\[3\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[1\]
+ _02882_ top_inst.grid_inst.data_path_wires\[17\]\[4\] VGND VGND VPWR VPWR _02944_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_160_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22183_ _03860_ _03872_ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21134_ _02885_ _02021_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21065_ net869 _01735_ _02829_ _02707_ VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20016_ _01827_ _01832_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_232_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_225_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21967_ top_inst.grid_inst.data_path_wires\[18\]\[0\] VGND VGND VPWR VPWR _03680_
+ sky130_fd_sc_hd__clkbuf_4
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23706_ clknet_leaf_124_clk _00239_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_20918_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[23\] _02470_ VGND
+ VGND VPWR VPWR _02688_ sky130_fd_sc_hd__nand2_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21898_ _03614_ _03615_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23637_ clknet_leaf_126_clk _00170_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20849_ _02596_ _02621_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14370_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _07074_ sky130_fd_sc_hd__buf_2
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23568_ clknet_leaf_103_clk _00101_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13321_ _05759_ _05757_ _05753_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22519_ _04137_ _04199_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23499_ clknet_leaf_141_clk _00032_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[89\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16040_ _08642_ _08644_ _08645_ _08647_ _05313_ VGND VGND VPWR VPWR _08648_ sky130_fd_sc_hd__o311a_1
XFILLER_0_107_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13252_ _05985_ _05982_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__and2b_1
XFILLER_0_161_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12203_ net768 _05129_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_889 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13183_ _05959_ _05961_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12134_ net506 _05084_ _05091_ _05088_ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__o211a_1
X_17991_ _10413_ _10493_ VGND VGND VPWR VPWR _10494_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19730_ _11177_ _01557_ _01558_ _11714_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16942_ _09489_ _09490_ VGND VGND VPWR VPWR _09497_ sky130_fd_sc_hd__nand2_1
X_12065_ net518 _05045_ _05052_ _05049_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_1072 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19661_ _01298_ _11695_ net194 top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_217_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16873_ _09361_ _09191_ net224 _09213_ VGND VGND VPWR VPWR _09430_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_204_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18612_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[14\] _10639_ VGND
+ VGND VPWR VPWR _11072_ sky130_fd_sc_hd__or2_1
XTAP_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15824_ _08143_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[7\] _08169_
+ _08163_ VGND VGND VPWR VPWR _08437_ sky130_fd_sc_hd__and4b_1
XFILLER_0_232_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19592_ _01392_ _01422_ _01423_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__nand3_1
XTAP_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ _10961_ _10962_ _10994_ VGND VGND VPWR VPWR _11004_ sky130_fd_sc_hd__a21o_1
X_12967_ _05738_ _05756_ _05760_ _05743_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__o211a_1
X_15755_ _08152_ _08150_ _08157_ _08155_ VGND VGND VPWR VPWR _08370_ sky130_fd_sc_hd__and4_1
XTAP_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14706_ _07392_ _07393_ _07363_ VGND VGND VPWR VPWR _07395_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_129_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _04874_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__clkbuf_4
X_18474_ _10935_ VGND VGND VPWR VPWR _10937_ sky130_fd_sc_hd__inv_2
X_12898_ _05298_ _05672_ _05702_ VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15686_ _08300_ _08301_ _08269_ VGND VGND VPWR VPWR _08303_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_185_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _09952_ _09962_ VGND VGND VPWR VPWR _09963_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14637_ _07289_ _07298_ VGND VGND VPWR VPWR _07327_ sky130_fd_sc_hd__and2_1
XFILLER_0_185_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11849_ _04874_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__buf_2
XFILLER_0_200_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17356_ _09625_ _09895_ VGND VGND VPWR VPWR _09897_ sky130_fd_sc_hd__nand2_1
X_14568_ _07213_ _07215_ VGND VGND VPWR VPWR _07260_ sky130_fd_sc_hd__and2b_1
XFILLER_0_166_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16307_ _08883_ _08888_ VGND VGND VPWR VPWR _08889_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13519_ _06267_ _06268_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__xor2_2
X_14499_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[1\] _07081_ _07085_
+ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _07192_ sky130_fd_sc_hd__a22o_1
X_17287_ _09822_ _09827_ VGND VGND VPWR VPWR _09831_ sky130_fd_sc_hd__or2b_1
X_19026_ _11402_ _11404_ _11403_ VGND VGND VPWR VPWR _11447_ sky130_fd_sc_hd__o21ba_1
X_16238_ _08792_ _08793_ _08820_ _08821_ VGND VGND VPWR VPWR _08822_ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16169_ _08749_ _08754_ VGND VGND VPWR VPWR _08755_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_228_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19928_ _01736_ _01748_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19859_ _01352_ _01353_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[17\]
+ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__or3b_1
XFILLER_0_236_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22870_ net728 _04517_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_1323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21821_ _03510_ _03523_ _03542_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24540_ clknet_leaf_102_clk _01073_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_148_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21752_ _03475_ _03476_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20703_ _02480_ _02481_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__or2b_1
X_24471_ clknet_leaf_37_clk _01004_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21683_ _03404_ _03410_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23422_ top_inst.axis_out_inst.out_buff_data\[100\] _04596_ VGND VGND VPWR VPWR _04832_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20634_ _02394_ _02414_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23353_ _04690_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20565_ top_inst.deskew_buff_inst.col_input\[42\] _11723_ _02346_ _02347_ VGND VGND
+ VPWR VPWR _02348_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22304_ _03987_ _03990_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_162_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23284_ _04690_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__clkbuf_4
X_20496_ _02278_ _02279_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22235_ _03877_ _03876_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__and2b_1
XFILLER_0_132_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22166_ _03851_ _03855_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21117_ top_inst.grid_inst.data_path_wires\[17\]\[5\] VGND VGND VPWR VPWR _02873_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22097_ _03690_ _03688_ _03700_ _03697_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__nand4_1
XFILLER_0_195_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21048_ _02643_ _02811_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__nor2_1
XFILLER_0_233_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13870_ _06602_ _06605_ _06540_ VGND VGND VPWR VPWR _06610_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12821_ _05591_ _05593_ _05628_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_9_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22999_ net903 _04588_ _04591_ _04590_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12752_ net1010 _05403_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__nand2_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15540_ _08163_ _07639_ _08165_ _08166_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__o211a_1
XFILLER_0_243_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15471_ _08110_ _08111_ VGND VGND VPWR VPWR _08112_ sky130_fd_sc_hd__xnor2_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _05492_ _05493_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _09752_ _09757_ VGND VGND VPWR VPWR _09758_ sky130_fd_sc_hd__xor2_2
X_14422_ _07105_ _07106_ _07108_ VGND VGND VPWR VPWR _07118_ sky130_fd_sc_hd__and3_1
XFILLER_0_182_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18190_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[3\] _05730_ VGND
+ VGND VPWR VPWR _10661_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14353_ top_inst.skew_buff_inst.row\[1\].output_reg\[0\] top_inst.axis_in_inst.inbuf_bus\[8\]
+ net206 VGND VGND VPWR VPWR _07060_ sky130_fd_sc_hd__mux2_4
X_17141_ _09690_ _09664_ VGND VGND VPWR VPWR _09692_ sky130_fd_sc_hd__or2b_1
XFILLER_0_128_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13304_ net1033 _05788_ _06079_ _05767_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__o211a_1
XFILLER_0_243_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17072_ _09623_ VGND VGND VPWR VPWR _09624_ sky130_fd_sc_hd__clkbuf_4
X_14284_ _05632_ _06994_ VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_243_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13235_ top_inst.grid_inst.data_path_wires\[1\]\[5\] _05768_ VGND VGND VPWR VPWR
+ _06012_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16023_ _08532_ _08630_ VGND VGND VPWR VPWR _08631_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13166_ _05759_ _05757_ top_inst.grid_inst.data_path_wires\[1\]\[7\] VGND VGND VPWR
+ VPWR _05945_ sky130_fd_sc_hd__o21ai_4
X_12117_ net510 _05071_ _05081_ _05075_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13097_ _05822_ _05876_ _05877_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__a21oi_1
X_17974_ _10408_ _10437_ _10435_ VGND VGND VPWR VPWR _10478_ sky130_fd_sc_hd__o21a_1
XFILLER_0_236_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19713_ _01539_ _01540_ _01488_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__o21ai_1
X_16925_ _09478_ _09479_ _09480_ VGND VGND VPWR VPWR _09481_ sky130_fd_sc_hd__nand3_2
X_12048_ net793 _05036_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__or2_1
XFILLER_0_236_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19644_ _01432_ _01466_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__or2_1
X_16856_ _09411_ _09412_ VGND VGND VPWR VPWR _09413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_204_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15807_ _08414_ _08420_ VGND VGND VPWR VPWR _08421_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_220_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19575_ _11701_ _11696_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__and2_1
XFILLER_0_215_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16787_ _09311_ _09344_ _09345_ VGND VGND VPWR VPWR _09346_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13999_ top_inst.grid_inst.data_path_wires\[3\]\[5\] top_inst.grid_inst.data_path_wires\[3\]\[4\]
+ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__and4_1
XFILLER_0_133_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18526_ _10933_ _10941_ _10987_ VGND VGND VPWR VPWR _10988_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_220_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15738_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _08353_ sky130_fd_sc_hd__inv_2
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18457_ _10071_ _10919_ _10920_ _10620_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__o211a_1
X_15669_ _08149_ top_inst.grid_inst.data_path_wires\[7\]\[5\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[1\]
+ _08154_ VGND VGND VPWR VPWR _08286_ sky130_fd_sc_hd__nand4_1
XFILLER_0_213_1083 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17408_ _09945_ _09946_ VGND VGND VPWR VPWR _09947_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18388_ _10595_ _10602_ VGND VGND VPWR VPWR _10853_ sky130_fd_sc_hd__nand2_4
XFILLER_0_185_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17339_ _09868_ _09879_ _09870_ VGND VGND VPWR VPWR _09881_ sky130_fd_sc_hd__nand3_1
XFILLER_0_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20350_ _01993_ _02015_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[6\]
+ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__nand3_1
XFILLER_0_125_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19009_ _11388_ _11392_ _11390_ VGND VGND VPWR VPWR _11430_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20281_ _02068_ _02069_ _02049_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_140_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22020_ _03715_ _03716_ _06178_ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23971_ clknet_leaf_86_clk _00504_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_215_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22922_ net732 _04543_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__or2_1
XFILLER_0_192_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22853_ net387 _04504_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_233_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_635 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21804_ _03311_ _03526_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22784_ _04451_ _04444_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__or2b_1
XFILLER_0_79_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24523_ clknet_leaf_128_clk _01056_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_213_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21735_ _03458_ _03459_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24454_ clknet_leaf_62_clk _00987_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21666_ _03339_ _03366_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_1319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23405_ net66 _04658_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20617_ _02003_ _02015_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[12\]
+ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__a21o_1
X_24385_ clknet_leaf_38_clk net716 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21597_ _03253_ _03327_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23336_ net159 _04779_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20548_ _02009_ VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23267_ net126 _04740_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__or2_1
X_20479_ _02221_ _02263_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13020_ _05792_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_1386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22218_ _03903_ _03906_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__xnor2_2
XTAP_6700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23198_ net93 _04701_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__or2_1
XTAP_6711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22149_ _03806_ _03838_ _03839_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__and3_1
XTAP_6744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14971_ _07610_ _06647_ _07632_ _07618_ VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__o211a_1
XFILLER_0_234_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16710_ _09268_ _09269_ _09267_ VGND VGND VPWR VPWR _09271_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_22_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13922_ _06648_ _06641_ VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17690_ _10198_ _10199_ VGND VGND VPWR VPWR _10200_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16641_ top_inst.skew_buff_inst.row\[2\].output_reg\[5\] top_inst.axis_in_inst.inbuf_bus\[21\]
+ _05265_ VGND VGND VPWR VPWR _09209_ sky130_fd_sc_hd__mux2_4
XFILLER_0_202_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13853_ _06562_ _06565_ _06592_ VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__and3_1
XFILLER_0_242_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12804_ _05573_ _05577_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__or2b_1
X_19360_ _01195_ _01196_ _01178_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__o21ai_1
X_16572_ _08831_ _09147_ VGND VGND VPWR VPWR _09148_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13784_ _06198_ _06212_ VGND VGND VPWR VPWR _06527_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18311_ _10737_ _10739_ VGND VGND VPWR VPWR _10778_ sky130_fd_sc_hd__nor2_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15523_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _08154_ sky130_fd_sc_hd__buf_2
X_12735_ _05542_ _05544_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__xor2_1
XFILLER_0_167_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19291_ net240 VGND VGND VPWR VPWR _11692_ sky130_fd_sc_hd__buf_4
XFILLER_0_123_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ _10710_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__clkbuf_1
X_12666_ _05476_ _05477_ _05435_ _05437_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__a211o_1
X_15454_ _08094_ _08095_ VGND VGND VPWR VPWR _08096_ sky130_fd_sc_hd__nand2_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14405_ net1045 _06660_ _07102_ _07092_ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18173_ _10577_ _10604_ _10602_ _10599_ VGND VGND VPWR VPWR _10644_ sky130_fd_sc_hd__a22o_1
X_12597_ _05389_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__inv_2
X_15385_ _08028_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17124_ _09213_ _09211_ _09219_ VGND VGND VPWR VPWR _09675_ sky130_fd_sc_hd__and3_1
XFILLER_0_167_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14336_ _07043_ _07044_ VGND VGND VPWR VPWR _07045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold508 top_inst.axis_out_inst.out_buff_data\[69\] VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__dlygate4sd3_1
X_17055_ _09604_ _09605_ _09606_ VGND VGND VPWR VPWR _09608_ sky130_fd_sc_hd__a21o_1
X_14267_ _06898_ net180 _06977_ VGND VGND VPWR VPWR _06978_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_122_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold519 _00094_ VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_243_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13218_ _05896_ _05898_ _05946_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__and3_1
X_16006_ _08580_ _08581_ VGND VGND VPWR VPWR _08615_ sky130_fd_sc_hd__or2b_1
X_14198_ _06865_ _06862_ VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__and2b_1
XFILLER_0_141_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13149_ top_inst.grid_inst.data_path_wires\[1\]\[2\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[6\]
+ _05926_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__and3_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _10037_ _10300_ _10459_ VGND VGND VPWR VPWR _10461_ sky130_fd_sc_hd__o21ai_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16908_ _09460_ _09463_ VGND VGND VPWR VPWR _09464_ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17888_ _10366_ _10393_ VGND VGND VPWR VPWR _10394_ sky130_fd_sc_hd__xor2_1
XFILLER_0_206_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19627_ _01440_ _01456_ _01457_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16839_ _09393_ _09394_ _09395_ VGND VGND VPWR VPWR _09397_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_221_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19558_ _01346_ _01381_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__or2b_4
XFILLER_0_221_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18509_ _10969_ _10970_ VGND VGND VPWR VPWR _10971_ sky130_fd_sc_hd__nor2_1
X_19489_ _01307_ _01321_ _01322_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__nand3_2
XFILLER_0_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21520_ _03252_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__buf_2
XFILLER_0_180_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21451_ _03130_ _03148_ _03185_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_90_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20402_ top_inst.grid_inst.data_path_wires\[16\]\[7\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[6\]
+ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _02188_ sky130_fd_sc_hd__and3_2
X_24170_ clknet_leaf_23_clk _00703_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21382_ _03101_ _03103_ VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23121_ net787 _04656_ _04661_ _04662_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__o211a_1
X_20333_ _02117_ _02118_ _02119_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__a21o_1
XFILLER_0_222_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23052_ net6 _04615_ _04622_ _04619_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20264_ _01992_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[1\] _02052_
+ _02053_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__and4_1
Xoutput39 net39 VGND VGND VPWR VPWR output_tdata[100] sky130_fd_sc_hd__clkbuf_4
XTAP_6007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22003_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _03705_ sky130_fd_sc_hd__buf_2
XTAP_6029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20195_ top_inst.grid_inst.data_path_wires\[16\]\[5\] VGND VGND VPWR VPWR _01999_
+ sky130_fd_sc_hd__buf_4
XTAP_5317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_892 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23954_ clknet_leaf_91_clk _00487_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22905_ top_inst.skew_buff_inst.row\[2\].output_reg\[0\] _04530_ VGND VGND VPWR VPWR
+ _04538_ sky130_fd_sc_hd__or2_1
XTAP_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23885_ clknet_leaf_64_clk _00418_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22836_ top_inst.skew_buff_inst.row\[3\].output_reg\[2\] _03691_ VGND VGND VPWR VPWR
+ _04499_ sky130_fd_sc_hd__or2_1
XFILLER_0_195_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_1092 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22767_ _04268_ _04395_ _04412_ _04415_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__o31a_1
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12520_ _05333_ _05334_ _05336_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__o21ai_1
X_24506_ clknet_leaf_128_clk _01039_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dfxtp_4
X_21718_ _03444_ VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__clkbuf_1
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22698_ _04092_ _04370_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _05270_ _05272_ _05277_ _05261_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__o211a_1
X_24437_ clknet_leaf_58_clk _00970_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_21649_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[16\] _03122_ VGND
+ VGND VPWR VPWR _03378_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15170_ _07818_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24368_ clknet_leaf_31_clk _00901_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[127\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12382_ net568 _05230_ _05232_ _05221_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__o211a_1
XANTENNA_90 net143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14121_ _06833_ _06835_ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__xnor2_2
X_23319_ net151 _04766_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_244_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_240_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24299_ clknet_leaf_138_clk _00832_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[74\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_238_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14052_ _05632_ _06768_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13003_ _05312_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__buf_8
XFILLER_0_197_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18860_ _11282_ _11283_ _11262_ VGND VGND VPWR VPWR _11285_ sky130_fd_sc_hd__a21oi_1
XTAP_6530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17811_ _10317_ _10318_ VGND VGND VPWR VPWR _10319_ sky130_fd_sc_hd__nor2_1
XTAP_6563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18791_ _11158_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[13\]\[1\]
+ top_inst.grid_inst.data_path_wires\[13\]\[0\] VGND VGND VPWR VPWR _11218_ sky130_fd_sc_hd__nand4_1
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17742_ _10025_ _10056_ _10212_ VGND VGND VPWR VPWR _10251_ sky130_fd_sc_hd__and3_1
XTAP_5873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14954_ _07619_ _07611_ _07620_ _07618_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__o211a_1
XTAP_5884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13905_ _06198_ _06634_ _06636_ _06446_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__o211a_1
XFILLER_0_216_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17673_ _10154_ _10155_ _10182_ _10183_ VGND VGND VPWR VPWR _10184_ sky130_fd_sc_hd__a211o_1
X_14885_ _07559_ _07568_ VGND VGND VPWR VPWR _07569_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19412_ _01245_ _01246_ _01218_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_72_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16624_ _09185_ _09192_ _09195_ _09184_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13836_ _06575_ _06577_ VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_1165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19343_ _01181_ VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16555_ _09126_ _09130_ VGND VGND VPWR VPWR _09131_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13767_ _06465_ _06469_ _06463_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_169_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15506_ _07610_ _06634_ _08141_ _08142_ VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__o211a_1
X_12718_ _05286_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19274_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _11678_ sky130_fd_sc_hd__buf_2
X_16486_ _09023_ _09022_ VGND VGND VPWR VPWR _09064_ sky130_fd_sc_hd__or2b_1
XFILLER_0_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13698_ _06409_ _06403_ _06442_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__nand3_1
XFILLER_0_155_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_890 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18225_ top_inst.grid_inst.data_path_wires\[12\]\[5\] top_inst.grid_inst.data_path_wires\[12\]\[4\]
+ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _10694_ sky130_fd_sc_hd__nand4_1
XFILLER_0_170_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15437_ _08005_ _08078_ VGND VGND VPWR VPWR _08079_ sky130_fd_sc_hd__nor2_1
X_12649_ _05446_ _05460_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18156_ _10577_ _10602_ VGND VGND VPWR VPWR _10628_ sky130_fd_sc_hd__nand2_1
X_15368_ _07969_ _07975_ _07968_ VGND VGND VPWR VPWR _08012_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17107_ _09621_ _09658_ VGND VGND VPWR VPWR _09659_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14319_ _06966_ _06998_ _06999_ VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__o21ba_1
Xhold305 _00153_ VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18087_ top_inst.grid_inst.data_path_wires\[12\]\[0\] VGND VGND VPWR VPWR _10577_
+ sky130_fd_sc_hd__clkbuf_4
Xhold316 _00107_ VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15299_ _07941_ _07943_ _05315_ VGND VGND VPWR VPWR _07945_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold327 _01169_ VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold338 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[9\] VGND
+ VGND VPWR VPWR net520 sky130_fd_sc_hd__dlygate4sd3_1
X_17038_ _09465_ _09550_ _09549_ VGND VGND VPWR VPWR _09591_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_180_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold349 top_inst.deskew_buff_inst.col_input\[98\] VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18989_ _11394_ _11395_ _11409_ VGND VGND VPWR VPWR _11411_ sky130_fd_sc_hd__and3_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20951_ _02473_ _02718_ _02719_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__and3_1
XFILLER_0_205_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23670_ clknet_leaf_116_clk net356 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20882_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[19\] _02559_ _02621_
+ _02619_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22621_ _04296_ _04297_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22552_ _04227_ _04230_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21503_ _03112_ _03157_ _03235_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22483_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[15\] _03937_ VGND
+ VGND VPWR VPWR _04165_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24222_ clknet_leaf_12_clk _00755_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21434_ top_inst.grid_inst.data_path_wires\[17\]\[6\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[17\]\[7\]
+ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24153_ clknet_leaf_18_clk _00686_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21365_ _03044_ _03056_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_110_clk clknet_4_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23104_ net653 _10541_ _04650_ _04643_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20316_ _02089_ _02102_ _02103_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24084_ clknet_leaf_87_clk _00617_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold850 top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[27\] VGND VGND
+ VPWR VPWR net1032 sky130_fd_sc_hd__dlygate4sd3_1
X_21296_ _02999_ _03004_ _03033_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__o21ai_1
Xhold861 top_inst.axis_in_inst.inbuf_bus\[28\] VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23035_ net30 _04601_ _04612_ _04606_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__o211a_1
Xhold872 top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[13\] VGND VGND
+ VPWR VPWR net1054 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold883 top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[12\] VGND VGND
+ VPWR VPWR net1065 sky130_fd_sc_hd__dlygate4sd3_1
X_20247_ _01989_ _01986_ _02011_ _02009_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__nand4_2
Xhold894 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[25\] VGND VGND
+ VPWR VPWR net1076 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20178_ _01986_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__clkbuf_4
XTAP_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23937_ clknet_leaf_80_clk _00470_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11951_ net733 _04977_ _04986_ _04981_ VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__o211a_1
XTAP_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ _07316_ _07354_ _07358_ _07314_ VGND VGND VPWR VPWR _07359_ sky130_fd_sc_hd__a22oi_4
XTAP_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11882_ net891 _04938_ _04947_ _04942_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23868_ clknet_leaf_78_clk _00401_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13621_ top_inst.grid_inst.data_path_wires\[2\]\[2\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[6\]
+ _06366_ VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22819_ _04466_ _04462_ _04474_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__a21o_1
X_23799_ clknet_leaf_70_clk _00332_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16340_ top_inst.grid_inst.data_path_wires\[8\]\[2\] top_inst.grid_inst.data_path_wires\[8\]\[3\]
+ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _08921_ sky130_fd_sc_hd__and4b_1
XFILLER_0_66_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13552_ _06190_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[2\] _06298_
+ _06299_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__nand4_1
XFILLER_0_27_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12503_ _05280_ _05279_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16271_ _08846_ _08853_ VGND VGND VPWR VPWR _08854_ sky130_fd_sc_hd__xnor2_1
X_13483_ _06219_ _06223_ _06232_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__or3_2
XFILLER_0_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18010_ _10476_ _10451_ VGND VGND VPWR VPWR _10513_ sky130_fd_sc_hd__and2b_1
X_15222_ _07858_ _07860_ VGND VGND VPWR VPWR _07869_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12434_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[30\] _05262_
+ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15153_ _07794_ _07801_ VGND VGND VPWR VPWR _07802_ sky130_fd_sc_hd__xnor2_1
X_12365_ net495 _05217_ _05223_ _05221_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_101_clk clknet_4_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14104_ _06817_ _06818_ VGND VGND VPWR VPWR _06819_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19961_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[22\] _01764_ VGND
+ VGND VPWR VPWR _01780_ sky130_fd_sc_hd__xnor2_2
X_15084_ _07732_ _07734_ VGND VGND VPWR VPWR _07735_ sky130_fd_sc_hd__xor2_1
XFILLER_0_240_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12296_ net858 _05178_ _05184_ _05182_ VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14035_ _06630_ _06640_ _06637_ top_inst.grid_inst.data_path_wires\[3\]\[6\] VGND
+ VGND VPWR VPWR _06752_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_129_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18912_ _11300_ _11306_ _11334_ VGND VGND VPWR VPWR _11335_ sky130_fd_sc_hd__a21o_1
XFILLER_0_201_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19892_ _01714_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_219_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18843_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[6\] _11267_ VGND
+ VGND VPWR VPWR _11268_ sky130_fd_sc_hd__xor2_2
XFILLER_0_235_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18774_ _11194_ _11201_ VGND VGND VPWR VPWR _11202_ sky130_fd_sc_hd__xnor2_1
XTAP_5670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15986_ _08152_ _08169_ _08167_ VGND VGND VPWR VPWR _08595_ sky130_fd_sc_hd__and3_1
XFILLER_0_234_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17725_ _10044_ _10042_ top_inst.grid_inst.data_path_wires\[11\]\[7\] VGND VGND VPWR
+ VPWR _10234_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14937_ top_inst.grid_inst.data_path_wires\[6\]\[1\] VGND VGND VPWR VPWR _07608_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17656_ _10127_ _10132_ VGND VGND VPWR VPWR _10167_ sky130_fd_sc_hd__or2b_1
X_14868_ _07550_ _07552_ VGND VGND VPWR VPWR _07553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16607_ _09165_ _09180_ VGND VGND VPWR VPWR _09181_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13819_ _06527_ _06560_ VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17587_ _10086_ _10079_ _10098_ VGND VGND VPWR VPWR _10101_ sky130_fd_sc_hd__and3_1
X_14799_ _07473_ VGND VGND VPWR VPWR _07485_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19326_ _11719_ _11720_ _08181_ VGND VGND VPWR VPWR _11721_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_169_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16538_ _09111_ _09113_ _09114_ VGND VGND VPWR VPWR _09115_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_161_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1025 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19257_ _11664_ _11670_ VGND VGND VPWR VPWR _11671_ sky130_fd_sc_hd__xnor2_1
X_16469_ _09045_ _09046_ VGND VGND VPWR VPWR _09047_ sky130_fd_sc_hd__xor2_1
XFILLER_0_116_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_1008 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18208_ _10675_ _10677_ VGND VGND VPWR VPWR _10678_ sky130_fd_sc_hd__xor2_2
XFILLER_0_72_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19188_ _11603_ _11604_ VGND VGND VPWR VPWR _11605_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_1236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18139_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _10614_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold102 top_inst.valid_pipe\[3\] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _00924_ VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold124 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[27\] VGND
+ VGND VPWR VPWR net306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold135 top_inst.axis_out_inst.out_buff_data\[13\] VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__dlygate4sd3_1
X_21150_ _02875_ _02881_ _02896_ _02880_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__o211a_1
Xhold146 _00132_ VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold157 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[30\] VGND
+ VGND VPWR VPWR net339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20101_ _01876_ _01913_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__nand2_1
Xhold168 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[19\] VGND
+ VGND VPWR VPWR net350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold179 _00013_ VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__dlygate4sd3_1
X_21081_ _02819_ _02843_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20032_ _01562_ _01846_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_238_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21983_ _06619_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__buf_4
XFILLER_0_197_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20934_ _02686_ _02703_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__xor2_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23722_ clknet_leaf_120_clk _00255_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23653_ clknet_leaf_128_clk net351 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_20865_ _06701_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_230_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22604_ _04253_ _04278_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23584_ clknet_leaf_106_clk net316 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20796_ _02541_ _02570_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22535_ _04163_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22466_ _04124_ _04125_ _04148_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21417_ _03121_ _03152_ VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__xnor2_1
X_24205_ clknet_leaf_117_clk _00738_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22397_ _04058_ _04081_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12150_ net686 _05089_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__or2_1
X_24136_ clknet_leaf_144_clk _00669_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21348_ _02873_ _02871_ _02891_ _02889_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__nand4_1
XFILLER_0_20_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24067_ clknet_leaf_84_clk _00600_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_12081_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[7\] _05050_
+ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold680 top_inst.deskew_buff_inst.col_input\[38\] VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__dlygate4sd3_1
X_21279_ _03006_ _03017_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_241_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold691 top_inst.axis_out_inst.out_buff_data\[53\] VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23018_ _04602_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15840_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[9\] _08452_ _08373_
+ VGND VGND VPWR VPWR _08453_ sky130_fd_sc_hd__a21o_1
XFILLER_0_244_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _08324_ _08331_ _08329_ VGND VGND VPWR VPWR _08386_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_231_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12983_ _05751_ _05756_ _05771_ _05767_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__o211a_1
XTAP_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ top_inst.grid_inst.data_path_wires\[11\]\[6\] VGND VGND VPWR VPWR _10037_
+ sky130_fd_sc_hd__buf_2
XTAP_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14722_ _07383_ _07384_ VGND VGND VPWR VPWR _07410_ sky130_fd_sc_hd__or2b_1
XTAP_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ net905 _04964_ _04976_ _04968_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__o211a_1
X_18490_ _10949_ _10951_ VGND VGND VPWR VPWR _10953_ sky130_fd_sc_hd__nand2_1
XTAP_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _09972_ _09977_ VGND VGND VPWR VPWR _09978_ sky130_fd_sc_hd__and2b_1
XFILLER_0_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14653_ _07326_ _07327_ _07341_ VGND VGND VPWR VPWR _07343_ sky130_fd_sc_hd__or3_1
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11865_ net897 _04925_ _04937_ _04929_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13604_ _06304_ _06312_ _06351_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__o21ai_1
X_17372_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[25\] _09631_ VGND
+ VGND VPWR VPWR _09912_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14584_ _07273_ _07274_ VGND VGND VPWR VPWR _07275_ sky130_fd_sc_hd__nand2_1
X_11796_ _04859_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19111_ _11479_ _11528_ VGND VGND VPWR VPWR _11530_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16323_ _08892_ _08904_ VGND VGND VPWR VPWR _08905_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13535_ _06259_ _06284_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__or2_1
X_19042_ _11427_ _11462_ VGND VGND VPWR VPWR _11463_ sky130_fd_sc_hd__nand2_1
X_16254_ _08835_ _08836_ VGND VGND VPWR VPWR _08837_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13466_ _06181_ _06202_ _06200_ _06184_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15205_ _07840_ _07852_ VGND VGND VPWR VPWR _07853_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12417_ net321 _05243_ _05252_ _05247_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16185_ _08764_ _08769_ VGND VGND VPWR VPWR _08770_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_211_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13397_ _06168_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__buf_8
XFILLER_0_112_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_1097 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15136_ _07783_ _07784_ VGND VGND VPWR VPWR _07785_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12348_ net879 _05204_ _05213_ _05208_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__o211a_1
X_19944_ _01480_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__buf_4
X_15067_ _07711_ _07716_ VGND VGND VPWR VPWR _07718_ sky130_fd_sc_hd__nand2_1
X_12279_ net691 _05169_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14018_ _06716_ _06719_ VGND VGND VPWR VPWR _06735_ sky130_fd_sc_hd__nand2_1
X_19875_ _01524_ _01683_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18826_ _11203_ _11224_ _11251_ VGND VGND VPWR VPWR _11252_ sky130_fd_sc_hd__o21ai_1
XTAP_6190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18757_ _11178_ _11184_ VGND VGND VPWR VPWR _11186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15969_ _08530_ _08537_ _08528_ VGND VGND VPWR VPWR _08579_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_234_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17708_ _10203_ _10217_ VGND VGND VPWR VPWR _10218_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18688_ _11132_ _11133_ VGND VGND VPWR VPWR _11134_ sky130_fd_sc_hd__or2_1
XFILLER_0_194_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_203_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17639_ _10125_ _10149_ _08265_ VGND VGND VPWR VPWR _10151_ sky130_fd_sc_hd__o21a_1
XFILLER_0_203_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20650_ _02004_ _02016_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[13\]
+ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__nand3_1
XFILLER_0_58_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19309_ _11703_ _05276_ _11706_ _11641_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20581_ _02355_ _02362_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22320_ _03887_ _03926_ _03972_ _04006_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22251_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[8\] _03937_ _03938_
+ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21202_ _02943_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22182_ _03865_ _03871_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21133_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _02885_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21064_ _02827_ _02828_ _06178_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20015_ _01831_ _01825_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__xor2_1
XFILLER_0_119_1200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_240_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_240_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21966_ net954 _03528_ _03677_ _03679_ _02962_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23705_ clknet_leaf_125_clk net529 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20917_ _02518_ _02668_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__and2_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21897_ _03279_ _03613_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20848_ _02619_ _02620_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__nor2_1
X_23636_ clknet_leaf_125_clk _00169_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23567_ clknet_leaf_103_clk _00100_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20779_ _02518_ _02554_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13320_ _06093_ _06094_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22518_ _04194_ _04198_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__xor2_1
XFILLER_0_162_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23498_ clknet_leaf_140_clk _00031_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[88\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13251_ _06023_ _06027_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22449_ _04127_ _04131_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12202_ net910 _05123_ _05130_ _05128_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13182_ _05911_ _05913_ _05960_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_20_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12133_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[29\] _05089_
+ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24119_ clknet_leaf_13_clk _00652_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_17990_ _10491_ _10492_ VGND VGND VPWR VPWR _10493_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16941_ _05326_ VGND VGND VPWR VPWR _09496_ sky130_fd_sc_hd__buf_8
X_12064_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[31\] _05050_
+ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19660_ _01297_ _01314_ _11695_ net235 VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__or4b_4
XFILLER_0_99_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16872_ _09360_ _09377_ _09191_ _09196_ VGND VGND VPWR VPWR _09429_ sky130_fd_sc_hd__or4b_4
X_18611_ _11040_ _11070_ VGND VGND VPWR VPWR _11071_ sky130_fd_sc_hd__xor2_1
XFILLER_0_189_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15823_ _08404_ _08410_ _08435_ VGND VGND VPWR VPWR _08436_ sky130_fd_sc_hd__o21a_1
XFILLER_0_176_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19591_ _01420_ _01421_ _01374_ _01393_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ _10952_ _10995_ _10996_ VGND VGND VPWR VPWR _11003_ sky130_fd_sc_hd__or3_1
XTAP_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15754_ _08366_ _08368_ VGND VGND VPWR VPWR _08369_ sky130_fd_sc_hd__xnor2_1
XTAP_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12966_ _05759_ _05294_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _07363_ _07392_ _07393_ VGND VGND VPWR VPWR _07394_ sky130_fd_sc_hd__and3_1
XTAP_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ net673 _04956_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18473_ _10934_ _10935_ _10592_ _10610_ VGND VGND VPWR VPWR _10936_ sky130_fd_sc_hd__and4b_1
XFILLER_0_157_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15685_ _08269_ _08300_ _08301_ VGND VGND VPWR VPWR _08302_ sky130_fd_sc_hd__and3_1
X_12897_ _05644_ _05673_ _05674_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__o21ba_1
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17424_ _09960_ _09961_ _09937_ VGND VGND VPWR VPWR _09962_ sky130_fd_sc_hd__mux2_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _07296_ _07297_ VGND VGND VPWR VPWR _07326_ sky130_fd_sc_hd__nor2_1
XFILLER_0_185_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11848_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[3\] _04917_
+ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _09624_ _09895_ VGND VGND VPWR VPWR _09896_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14567_ _07256_ _07257_ net230 _07198_ VGND VGND VPWR VPWR _07259_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11779_ _04874_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__buf_2
XFILLER_0_138_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16306_ _08886_ _08887_ VGND VGND VPWR VPWR _08888_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13518_ top_inst.grid_inst.data_path_wires\[2\]\[3\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[2\]
+ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__and2_1
X_17286_ _09807_ _09821_ VGND VGND VPWR VPWR _09830_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14498_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[5\] _07163_ _07164_
+ VGND VGND VPWR VPWR _07191_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_126_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19025_ _11442_ _11445_ VGND VGND VPWR VPWR _11446_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16237_ _08818_ _08819_ _08794_ _08795_ VGND VGND VPWR VPWR _08821_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13449_ _06208_ _05773_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16168_ _08750_ _08753_ VGND VGND VPWR VPWR _08754_ sky130_fd_sc_hd__xor2_2
XFILLER_0_23_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15119_ _07743_ _07744_ _07767_ _07768_ VGND VGND VPWR VPWR _07769_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_228_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16099_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _08693_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19927_ _01746_ _01747_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_227_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19858_ _01524_ _01659_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18809_ _11233_ _11234_ VGND VGND VPWR VPWR _11235_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_1302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19789_ _01614_ _01615_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21820_ _03519_ _03541_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21751_ _03278_ _03474_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_90_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20702_ _02479_ _02477_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__or2b_1
X_24470_ clknet_leaf_55_clk _01003_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_21682_ _03405_ _03409_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23421_ net318 _04827_ _04830_ _04831_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__o211a_1
X_20633_ _02411_ _02413_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_4_9__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_4_9__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23352_ net40 _04792_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20564_ _02343_ _02345_ _10831_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22303_ _03988_ _03989_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_190_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23283_ net134 _04753_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20495_ _01993_ _02229_ _02276_ _02277_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__nor4_1
XFILLER_0_132_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22234_ _03919_ _03922_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22165_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[7\] _03854_ VGND
+ VGND VPWR VPWR _03855_ sky130_fd_sc_hd__xor2_2
XFILLER_0_203_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21116_ _01997_ _11142_ _02872_ _02707_ VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__o211a_1
X_22096_ top_inst.grid_inst.data_path_wires\[18\]\[4\] top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[1\]
+ _03697_ _03690_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__a22o_1
XFILLER_0_227_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21047_ _02643_ _02811_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12820_ _05626_ _05627_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_198_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22998_ top_inst.skew_buff_inst.row\[0\].output_reg\[0\] _04583_ VGND VGND VPWR VPWR
+ _04591_ sky130_fd_sc_hd__or2_1
XFILLER_0_241_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ net1084 _05314_ _05560_ _05308_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__o211a_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21949_ _03549_ _03643_ _03645_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_243_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_81_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15470_ _08077_ _08080_ _08079_ VGND VGND VPWR VPWR _08111_ sky130_fd_sc_hd__o21ba_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12682_ _05298_ _05287_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__nand2_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14421_ _04869_ VGND VGND VPWR VPWR _07117_ sky130_fd_sc_hd__clkbuf_4
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23619_ clknet_leaf_102_clk net502 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24599_ clknet_leaf_23_clk _01132_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_33_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17140_ _09664_ _09690_ VGND VGND VPWR VPWR _09691_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14352_ net34 VGND VGND VPWR VPWR _07059_ sky130_fd_sc_hd__buf_8
XFILLER_0_170_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_971 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13303_ _06077_ _06078_ _05328_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__a21o_1
X_17071_ _09591_ VGND VGND VPWR VPWR _09623_ sky130_fd_sc_hd__buf_4
X_14283_ _06960_ _06993_ _05316_ VGND VGND VPWR VPWR _06994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16022_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[15\] _08452_ VGND
+ VGND VPWR VPWR _08630_ sky130_fd_sc_hd__xnor2_2
X_13234_ _06009_ _06010_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13165_ _05751_ _05904_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12116_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[22\] _05076_
+ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__or2_1
X_13096_ _05839_ _05838_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__and2b_1
X_17973_ _10451_ _10476_ VGND VGND VPWR VPWR _10477_ sky130_fd_sc_hd__xor2_1
XFILLER_0_209_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16924_ _09427_ _09435_ _09434_ VGND VGND VPWR VPWR _09480_ sky130_fd_sc_hd__a21bo_1
X_19712_ _01488_ _01539_ _01540_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__or3_1
XFILLER_0_40_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12047_ net696 _05031_ _05041_ _05035_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__o211a_1
XFILLER_0_237_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16855_ _09362_ _09368_ VGND VGND VPWR VPWR _09412_ sky130_fd_sc_hd__or2b_1
X_19643_ _01473_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_233_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15806_ _08415_ _08419_ VGND VGND VPWR VPWR _08420_ sky130_fd_sc_hd__xor2_1
XFILLER_0_88_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19574_ _01402_ _01405_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__xor2_2
X_16786_ _09331_ _09332_ _09342_ _09343_ VGND VGND VPWR VPWR _09345_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13998_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[2\] _06624_ _06693_
+ _06692_ top_inst.grid_inst.data_path_wires\[3\]\[0\] VGND VGND VPWR VPWR _06716_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18525_ _10936_ _10938_ _10940_ VGND VGND VPWR VPWR _10987_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15737_ top_inst.grid_inst.data_path_wires\[7\]\[1\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[7\]
+ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[7\]\[2\]
+ VGND VGND VPWR VPWR _08352_ sky130_fd_sc_hd__and4b_1
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12949_ _05746_ _05735_ _05747_ _05743_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__o211a_1
XFILLER_0_220_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18456_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[10\] _10639_ VGND
+ VGND VPWR VPWR _10920_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15668_ top_inst.grid_inst.data_path_wires\[7\]\[5\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[1\]
+ _08154_ top_inst.grid_inst.data_path_wires\[7\]\[6\] VGND VGND VPWR VPWR _08285_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17407_ _09933_ _09944_ VGND VGND VPWR VPWR _09946_ sky130_fd_sc_hd__nand2_1
Xclkbuf_2_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_14619_ _07308_ _07309_ VGND VGND VPWR VPWR _07310_ sky130_fd_sc_hd__and2_1
XFILLER_0_185_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18387_ _10849_ _10851_ VGND VGND VPWR VPWR _10852_ sky130_fd_sc_hd__and2_1
X_15599_ _08218_ VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17338_ _09868_ _09870_ _09879_ VGND VGND VPWR VPWR _09880_ sky130_fd_sc_hd__a21o_1
XFILLER_0_185_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17269_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[20\] _09631_ VGND
+ VGND VPWR VPWR _09814_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_1150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19008_ _11416_ _11386_ VGND VGND VPWR VPWR _11429_ sky130_fd_sc_hd__or2b_1
XFILLER_0_125_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20280_ _02049_ _02068_ _02069_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_209_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23970_ clknet_leaf_85_clk _00503_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_194_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22921_ net712 _04535_ _04546_ _04537_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22852_ net942 _04496_ _04507_ _04498_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_211_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21803_ top_inst.deskew_buff_inst.col_input\[86\] _05731_ _03510_ _03525_ VGND VGND
+ VPWR VPWR _03526_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22783_ _04444_ _04451_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__or2b_1
XFILLER_0_190_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_63_clk clknet_4_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24522_ clknet_leaf_131_clk _01055_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dfxtp_4
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21734_ _03458_ _03459_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__nor2_1
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24453_ clknet_leaf_62_clk _00986_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_21665_ _03392_ _03393_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23404_ net801 _04655_ _04822_ _04819_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20616_ _02004_ _02016_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[12\]
+ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__nand3_1
X_24384_ clknet_leaf_39_clk _00917_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21596_ _02897_ _02895_ _02878_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23335_ net831 _04778_ _04784_ _04782_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__o211a_1
X_20547_ _02328_ _02329_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23266_ net1023 _04739_ _04745_ _04743_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__o211a_1
X_20478_ _02262_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22217_ _03904_ _03905_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23197_ net673 _04700_ _04706_ _04704_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22148_ _03836_ _03837_ _03807_ _03808_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__o211ai_1
XTAP_6734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14970_ _07631_ _07075_ VGND VGND VPWR VPWR _07632_ sky130_fd_sc_hd__or2_1
X_22079_ _03771_ _03740_ _03749_ _03748_ _03747_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_233_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13921_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _06648_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16640_ _09185_ _09206_ _09208_ _09184_ VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13852_ _06562_ _06565_ _06592_ VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_230_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12803_ _05609_ _05610_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16571_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[14\] _08066_ _09145_
+ _09146_ VGND VGND VPWR VPWR _09147_ sky130_fd_sc_hd__a22o_1
X_13783_ _06193_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[7\] _06214_
+ _06195_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__and4b_1
XFILLER_0_198_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_54_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18310_ _10751_ _10776_ VGND VGND VPWR VPWR _10777_ sky130_fd_sc_hd__xnor2_1
X_15522_ _07624_ _06634_ _08153_ _08142_ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__o211a_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19290_ top_inst.skew_buff_inst.row\[3\].output_reg\[3\] top_inst.axis_in_inst.inbuf_bus\[27\]
+ net184 VGND VGND VPWR VPWR _11691_ sky130_fd_sc_hd__mux2_4
X_12734_ _05496_ _05501_ _05543_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18241_ _10641_ _10709_ VGND VGND VPWR VPWR _10710_ sky130_fd_sc_hd__and2_1
X_15453_ _08016_ _08018_ _08060_ _08061_ _08063_ VGND VGND VPWR VPWR _08095_ sky130_fd_sc_hd__a32o_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12665_ _05474_ _05475_ _05441_ _05442_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__a211o_1
XFILLER_0_132_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14404_ _07100_ _07101_ _05336_ VGND VGND VPWR VPWR _07102_ sky130_fd_sc_hd__o21ai_1
X_18172_ _10632_ _10633_ VGND VGND VPWR VPWR _10643_ sky130_fd_sc_hd__or2b_1
XFILLER_0_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15384_ _07117_ _08027_ VGND VGND VPWR VPWR _08028_ sky130_fd_sc_hd__and2_1
X_12596_ _05391_ _05393_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17123_ _09597_ _09637_ _09636_ VGND VGND VPWR VPWR _09674_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_142_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14335_ _07020_ _07021_ _07018_ VGND VGND VPWR VPWR _07044_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_68_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17054_ _09604_ _09605_ _09606_ VGND VGND VPWR VPWR _09607_ sky130_fd_sc_hd__nand3_1
XFILLER_0_68_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold509 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[28\] VGND
+ VGND VPWR VPWR net691 sky130_fd_sc_hd__dlygate4sd3_1
X_14266_ _06640_ _06637_ _06635_ VGND VGND VPWR VPWR _06977_ sky130_fd_sc_hd__o21a_1
XFILLER_0_243_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16005_ _08612_ _08613_ VGND VGND VPWR VPWR _08614_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_106_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13217_ _05992_ _05994_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14197_ _06905_ _06909_ VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _05741_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[6\] _05926_
+ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__a21oi_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13079_ _05746_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[2\] _05857_
+ _05858_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__nand4_1
X_17956_ _10037_ _10300_ _10459_ VGND VGND VPWR VPWR _10460_ sky130_fd_sc_hd__or3_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16907_ _09461_ _09462_ VGND VGND VPWR VPWR _09463_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17887_ _10391_ _10392_ VGND VGND VPWR VPWR _10393_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19626_ _01453_ _01454_ _01455_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__a21o_1
X_16838_ _09393_ _09394_ _09395_ VGND VGND VPWR VPWR _09396_ sky130_fd_sc_hd__nor3_2
XFILLER_0_233_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16769_ _09325_ _09326_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[6\]
+ VGND VGND VPWR VPWR _09328_ sky130_fd_sc_hd__a21oi_1
X_19557_ _01345_ _01384_ _01388_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_177_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_45_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_221_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18508_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[12\] _10793_ VGND
+ VGND VPWR VPWR _10970_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19488_ _01319_ _01320_ _01312_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_927 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18439_ _10895_ _10902_ VGND VGND VPWR VPWR _10903_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21450_ _03145_ _03147_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__and2b_1
XFILLER_0_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20401_ _01989_ _02020_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21381_ _03105_ _03108_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__or2_2
XFILLER_0_86_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23120_ _04550_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__clkbuf_4
X_20332_ _02117_ _02118_ _02119_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__nand3_2
XFILLER_0_226_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23051_ net583 _04616_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20263_ top_inst.grid_inst.data_path_wires\[16\]\[0\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[3\]
+ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[2\] top_inst.grid_inst.data_path_wires\[16\]\[1\]
+ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22002_ _03684_ _05270_ _03704_ _03702_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__o211a_1
XTAP_6019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20194_ _01997_ _10033_ _01998_ _01840_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__o211a_1
XTAP_5307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23953_ clknet_leaf_90_clk _00486_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_231_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22904_ net764 _04535_ _04536_ _04537_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__o211a_1
XTAP_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23884_ clknet_leaf_61_clk _00417_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22835_ net578 _04496_ _04497_ _04498_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_233_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_36_clk clknet_4_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22766_ _04434_ _04435_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__or2_1
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24505_ clknet_leaf_126_clk _01038_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfxtp_4
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21717_ _03311_ _03443_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__and2_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22697_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[24\] _04163_ VGND
+ VGND VPWR VPWR _04370_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24436_ clknet_leaf_54_clk _00969_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12450_ _05273_ _05276_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21648_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[15\] _03376_ _03123_
+ VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24367_ clknet_leaf_31_clk _00900_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[126\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12381_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[8\] _05222_
+ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_80 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21579_ _03070_ _03309_ _03310_ _02909_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_91 net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14120_ _06782_ _06791_ _06834_ VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23318_ net658 _04765_ _04774_ _04769_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24298_ clknet_leaf_137_clk _00831_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14051_ _06734_ _06765_ _06766_ _06767_ VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__o31a_1
X_23249_ net838 _04726_ _04735_ _04730_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13002_ net1087 _05314_ _05786_ _05767_ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__o211a_1
XTAP_6520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17810_ _10314_ _10316_ VGND VGND VPWR VPWR _10318_ sky130_fd_sc_hd__and2_1
XTAP_6564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18790_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[2\] _11135_ VGND
+ VGND VPWR VPWR _11217_ sky130_fd_sc_hd__nand2_2
XFILLER_0_98_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17741_ _10245_ _10249_ VGND VGND VPWR VPWR _10250_ sky130_fd_sc_hd__xnor2_1
XTAP_5863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14953_ _04865_ _07416_ VGND VGND VPWR VPWR _07620_ sky130_fd_sc_hd__nand2_1
XTAP_5874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13904_ _06635_ _06620_ VGND VGND VPWR VPWR _06636_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17672_ _10180_ _10181_ _10156_ _10157_ VGND VGND VPWR VPWR _10183_ sky130_fd_sc_hd__o211a_1
X_14884_ _07566_ _07567_ VGND VGND VPWR VPWR _07568_ sky130_fd_sc_hd__nor2_1
XFILLER_0_215_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16623_ _09194_ _08684_ VGND VGND VPWR VPWR _09195_ sky130_fd_sc_hd__or2_1
X_19411_ _01245_ _01246_ _01218_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13835_ _06507_ _06545_ _06576_ VGND VGND VPWR VPWR _06577_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_clk clknet_4_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_187_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16554_ _09128_ _09129_ VGND VGND VPWR VPWR _09130_ sky130_fd_sc_hd__nor2_1
X_19342_ _11722_ _01180_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__and2_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13766_ _06505_ _06509_ VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_174_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15505_ _07617_ VGND VGND VPWR VPWR _08142_ sky130_fd_sc_hd__clkbuf_4
X_12717_ _05304_ _05490_ _05287_ _05302_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__a22o_1
X_19273_ net245 VGND VGND VPWR VPWR _11677_ sky130_fd_sc_hd__buf_2
X_16485_ _09061_ _09062_ VGND VGND VPWR VPWR _09063_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13697_ _06409_ _06403_ _06442_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18224_ top_inst.grid_inst.data_path_wires\[12\]\[4\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[12\]\[5\]
+ VGND VGND VPWR VPWR _10693_ sky130_fd_sc_hd__a22o_1
X_15436_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[14\] _07924_ VGND
+ VGND VPWR VPWR _08078_ sky130_fd_sc_hd__xnor2_1
X_12648_ _05454_ _05459_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__xor2_1
XFILLER_0_170_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18155_ net935 _10616_ _10627_ _10620_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__o211a_1
XFILLER_0_182_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15367_ _08003_ _08010_ VGND VGND VPWR VPWR _08011_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12579_ _05339_ _05360_ _05392_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__a21o_1
XFILLER_0_182_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17106_ _09622_ _09657_ VGND VGND VPWR VPWR _09658_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14318_ _06635_ _06652_ _06650_ VGND VGND VPWR VPWR _07027_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18086_ net646 _10563_ _10576_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__o21a_1
X_15298_ _07941_ _07943_ VGND VGND VPWR VPWR _07944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold306 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[10\] VGND
+ VGND VPWR VPWR net488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 top_inst.deskew_buff_inst.col_input\[127\] VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[22\] VGND
+ VGND VPWR VPWR net510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17037_ _09588_ _09589_ VGND VGND VPWR VPWR _09590_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold339 _00080_ VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__dlygate4sd3_1
X_14249_ net1090 VGND VGND VPWR VPWR _06960_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _11394_ _11395_ _11409_ VGND VGND VPWR VPWR _11410_ sky130_fd_sc_hd__a21oi_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _10404_ _10442_ VGND VGND VPWR VPWR _10444_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20950_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[24\] _02468_ VGND
+ VGND VPWR VPWR _02719_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19609_ _01436_ _01439_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__xor2_1
XFILLER_0_221_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20881_ _02651_ _02652_ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__and2_1
XFILLER_0_191_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_clk clknet_4_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22620_ _04271_ _04295_ _04286_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__nand3_1
XFILLER_0_221_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22551_ _04227_ _04230_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21502_ _03190_ _03231_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__and2_1
X_22482_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[14\] _04163_ _03938_
+ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__a21o_1
XFILLER_0_228_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24221_ clknet_leaf_118_clk _00754_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21433_ top_inst.grid_inst.data_path_wires\[17\]\[7\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _03168_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24152_ clknet_leaf_18_clk _00685_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_21364_ _03083_ _03100_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_130_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23103_ net354 _05323_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__or2_1
X_20315_ _01990_ _02016_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[5\]
+ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21295_ _02998_ _03005_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__or2b_1
X_24083_ clknet_leaf_87_clk _00616_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold840 top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[17\] VGND VGND
+ VPWR VPWR net1022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold851 top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[11\] VGND VGND
+ VPWR VPWR net1033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[0\] VGND VGND
+ VPWR VPWR net1044 sky130_fd_sc_hd__dlygate4sd3_1
X_23034_ net1112 _04603_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__or2_1
Xhold873 top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[15\] VGND VGND
+ VPWR VPWR net1055 sky130_fd_sc_hd__dlygate4sd3_1
X_20246_ _01986_ _02011_ _02009_ _01989_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__a22o_1
XFILLER_0_229_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold884 top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[13\] VGND VGND
+ VPWR VPWR net1066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold895 top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[0\] VGND VGND
+ VPWR VPWR net1077 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20177_ top_inst.grid_inst.data_path_wires\[16\]\[0\] VGND VGND VPWR VPWR _01986_
+ sky130_fd_sc_hd__buf_2
XTAP_5126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23936_ clknet_leaf_80_clk _00469_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ net651 _04982_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1057 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_1420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23867_ clknet_leaf_78_clk _00400_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11881_ net576 _04943_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13620_ _06186_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[6\] _06366_
+ VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__a21oi_1
X_22818_ _04449_ _04469_ _04482_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23798_ clknet_leaf_70_clk _00331_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_211_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13551_ _06190_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[2\] _06298_
+ _06299_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22749_ _04401_ _04419_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12502_ _05280_ _05272_ _05279_ _05273_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__a22o_1
X_16270_ _08851_ _08852_ VGND VGND VPWR VPWR _08853_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13482_ _06186_ _06202_ _06200_ _06188_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15221_ _07820_ _07864_ _07862_ VGND VGND VPWR VPWR _07868_ sky130_fd_sc_hd__a21bo_1
X_24419_ clknet_leaf_55_clk net663 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12433_ _05142_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__buf_4
XFILLER_0_81_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15152_ _07799_ _07800_ VGND VGND VPWR VPWR _07801_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12364_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[0\] _05222_
+ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14103_ _06632_ _06643_ _06815_ _06816_ VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__and4_1
XFILLER_0_239_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19960_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[21\] _01761_ _01762_
+ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__a21o_1
X_15083_ _07681_ _07703_ _07733_ VGND VGND VPWR VPWR _07734_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12295_ net848 _05183_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14034_ top_inst.grid_inst.data_path_wires\[3\]\[6\] top_inst.grid_inst.data_path_wires\[3\]\[5\]
+ _06640_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _06751_ sky130_fd_sc_hd__and4_2
X_18911_ _11301_ _11305_ VGND VGND VPWR VPWR _11334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_1408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19891_ _11722_ _01713_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18842_ _11265_ _11266_ VGND VGND VPWR VPWR _11267_ sky130_fd_sc_hd__nand2_1
XTAP_6350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18773_ _11199_ _11200_ VGND VGND VPWR VPWR _11201_ sky130_fd_sc_hd__xnor2_2
X_15985_ _08563_ _08562_ VGND VGND VPWR VPWR _08594_ sky130_fd_sc_hd__or2b_1
XFILLER_0_209_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14936_ _07606_ _05735_ _07607_ _07092_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__o211a_1
X_17724_ _10206_ _10208_ VGND VGND VPWR VPWR _10233_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14867_ _07444_ _07479_ _07517_ _07551_ VGND VGND VPWR VPWR _07552_ sky130_fd_sc_hd__a31o_1
XFILLER_0_199_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17655_ _10159_ _10165_ VGND VGND VPWR VPWR _10166_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16606_ _09174_ _09179_ VGND VGND VPWR VPWR _09180_ sky130_fd_sc_hd__xnor2_1
X_13818_ _06558_ _06559_ VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__nor2_1
X_17586_ _10099_ VGND VGND VPWR VPWR _10100_ sky130_fd_sc_hd__inv_2
X_14798_ _07477_ _07446_ VGND VGND VPWR VPWR _07484_ sky130_fd_sc_hd__or2b_4
XFILLER_0_169_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16537_ _09111_ _09113_ _05406_ VGND VGND VPWR VPWR _09114_ sky130_fd_sc_hd__a21oi_1
X_19325_ _11717_ _11718_ _11712_ VGND VGND VPWR VPWR _11720_ sky130_fd_sc_hd__nor3b_1
X_13749_ _06210_ _06208_ _06198_ VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19256_ _11666_ _11669_ VGND VGND VPWR VPWR _11670_ sky130_fd_sc_hd__xnor2_1
X_16468_ _08677_ _08695_ _09009_ _09008_ VGND VGND VPWR VPWR _09046_ sky130_fd_sc_hd__a31o_1
XFILLER_0_183_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15419_ _07982_ _08021_ VGND VGND VPWR VPWR _08062_ sky130_fd_sc_hd__and2b_1
X_18207_ _10652_ _10653_ _10676_ VGND VGND VPWR VPWR _10677_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_186_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19187_ _11563_ _11566_ _11602_ VGND VGND VPWR VPWR _11604_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16399_ _08977_ _08978_ VGND VGND VPWR VPWR _08979_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18138_ _10592_ _10607_ _10613_ _10594_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__o211a_1
XFILLER_0_182_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold103 _01019_ VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold114 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[3\] VGND VGND
+ VPWR VPWR net296 sky130_fd_sc_hd__dlygate4sd3_1
X_18069_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[16\] _10283_ _10234_
+ VGND VGND VPWR VPWR _10569_ sky130_fd_sc_hd__o21ba_1
Xhold125 _00258_ VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold136 top_inst.deskew_buff_inst.col_input\[99\] VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_7_clk clknet_4_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_223_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold147 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[19\] VGND
+ VGND VPWR VPWR net329 sky130_fd_sc_hd__dlygate4sd3_1
X_20100_ _01783_ _01896_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__nor2_1
Xhold158 _00197_ VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold169 _00186_ VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__dlygate4sd3_1
X_21080_ _02815_ _02842_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__xor2_1
XFILLER_0_229_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20031_ _01561_ _01846_ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_226_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21982_ top_inst.grid_inst.data_path_wires\[18\]\[5\] VGND VGND VPWR VPWR _03690_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23721_ clknet_leaf_121_clk _00254_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20933_ _02678_ _02702_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23652_ clknet_leaf_128_clk net342 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20864_ _02632_ _02636_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22603_ net542 _03528_ _04279_ _04280_ _09806_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__o221a_1
XFILLER_0_49_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23583_ clknet_leaf_110_clk _00116_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20795_ _02535_ _02565_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__or2b_1
XFILLER_0_130_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_863 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22534_ _04194_ _04198_ _04196_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22465_ _04126_ _04147_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24204_ clknet_leaf_16_clk _00737_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_888 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21416_ _03149_ _03151_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22396_ _04079_ _04080_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_241_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24135_ clknet_leaf_144_clk _00668_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21347_ _02871_ _02891_ _02889_ _02873_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24066_ clknet_leaf_84_clk _00599_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12080_ net458 _05058_ _05060_ _05049_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__o211a_1
Xhold670 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[0\] VGND VGND
+ VPWR VPWR net852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21278_ _03007_ _03016_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__xor2_1
Xhold681 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[19\] VGND
+ VGND VPWR VPWR net863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[5\] VGND
+ VGND VPWR VPWR net874 sky130_fd_sc_hd__dlygate4sd3_1
X_23017_ net33 net37 VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__and2_1
X_20229_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[7\] _02021_ VGND
+ VGND VPWR VPWR _02023_ sky130_fd_sc_hd__or2_1
XFILLER_0_200_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_232_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15770_ _08382_ _08384_ VGND VGND VPWR VPWR _08385_ sky130_fd_sc_hd__xnor2_1
X_12982_ _05770_ _05294_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__or2_1
XTAP_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _07405_ _07408_ VGND VGND VPWR VPWR _07409_ sky130_fd_sc_hd__xnor2_1
XTAP_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23919_ clknet_leaf_77_clk _00452_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ net595 _04969_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__or2_1
XTAP_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17440_ _09958_ _09976_ VGND VGND VPWR VPWR _09977_ sky130_fd_sc_hd__xnor2_1
XTAP_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14652_ _07326_ _07327_ _07341_ VGND VGND VPWR VPWR _07342_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_196_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11864_ net866 _04930_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__or2_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _06294_ _06303_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__or2_1
X_17371_ _09894_ _09897_ _09896_ VGND VGND VPWR VPWR _09911_ sky130_fd_sc_hd__a21o_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14583_ _07227_ _07233_ VGND VGND VPWR VPWR _07274_ sky130_fd_sc_hd__or2b_1
XFILLER_0_89_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11795_ net857 _04885_ _04897_ _04889_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16322_ _08902_ _08903_ VGND VGND VPWR VPWR _08904_ sky130_fd_sc_hd__nor2_1
X_19110_ _11479_ _11528_ VGND VGND VPWR VPWR _11529_ sky130_fd_sc_hd__nand2_1
X_13534_ _06281_ _06283_ VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19041_ _11460_ _11461_ VGND VGND VPWR VPWR _11462_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16253_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[5\] top_inst.grid_inst.data_path_wires\[8\]\[2\]
+ VGND VGND VPWR VPWR _08836_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13465_ _06184_ _06202_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15204_ _07850_ _07851_ VGND VGND VPWR VPWR _07852_ sky130_fd_sc_hd__nor2_1
X_12416_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[23\] _05248_
+ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__or2_1
X_16184_ _08767_ _08768_ VGND VGND VPWR VPWR _08769_ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13396_ _05312_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__buf_8
XFILLER_0_140_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15135_ top_inst.grid_inst.data_path_wires\[6\]\[2\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[5\]
+ VGND VGND VPWR VPWR _07784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12347_ net276 _05209_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19943_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[20\] _01761_ _01762_
+ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__a21o_1
X_15066_ _07711_ _07716_ VGND VGND VPWR VPWR _07717_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12278_ net981 _05164_ _05173_ _05168_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__o211a_1
X_14017_ _05633_ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__buf_8
XFILLER_0_142_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19874_ _01682_ _01687_ _01685_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_219_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18825_ _11222_ _11223_ VGND VGND VPWR VPWR _11251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_235_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18756_ _11178_ _11184_ VGND VGND VPWR VPWR _11185_ sky130_fd_sc_hd__or2_1
XTAP_5490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15968_ _08576_ _08577_ VGND VGND VPWR VPWR _08578_ sky130_fd_sc_hd__nor2_1
X_17707_ _10204_ _10216_ VGND VGND VPWR VPWR _10217_ sky130_fd_sc_hd__xnor2_1
X_14919_ net229 _07598_ _07594_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15899_ _08509_ _08510_ VGND VGND VPWR VPWR _08511_ sky130_fd_sc_hd__and2_1
X_18687_ _06619_ VGND VGND VPWR VPWR _11133_ sky130_fd_sc_hd__buf_2
XFILLER_0_76_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_203_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17638_ _10125_ _10149_ VGND VGND VPWR VPWR _10150_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17569_ _10083_ _05403_ VGND VGND VPWR VPWR _10084_ sky130_fd_sc_hd__nand2_1
XFILLER_0_175_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19308_ _05269_ _11705_ VGND VGND VPWR VPWR _11706_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20580_ _02356_ _02361_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19239_ _11624_ _11627_ _11652_ VGND VGND VPWR VPWR _11654_ sky130_fd_sc_hd__or3_1
XFILLER_0_144_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22250_ _03891_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21201_ _02135_ _02942_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__and2_1
XFILLER_0_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22181_ _03823_ _03870_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21132_ _02862_ _02881_ _02884_ _02880_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1086 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21063_ _02807_ _02809_ _02826_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__and3_1
X_20014_ _01828_ _01830_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__xor2_2
XFILLER_0_198_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21965_ _06178_ _03678_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__nand2_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23704_ clknet_leaf_125_clk net555 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ _02685_ _02664_ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__or2b_1
XFILLER_0_179_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21896_ _03279_ _03613_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_221_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23635_ clknet_leaf_108_clk net433 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_20847_ _02617_ _02618_ _02473_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23566_ clknet_leaf_103_clk net552 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20778_ _02520_ _02553_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22517_ _04196_ _04197_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23497_ clknet_leaf_142_clk _00030_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[87\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13250_ _06025_ _06026_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22448_ _04129_ _04130_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__and2b_1
XFILLER_0_17_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12201_ net723 _05129_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13181_ _05914_ _05915_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__or2b_1
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22379_ _04059_ _04063_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12132_ net266 _05084_ _05090_ _05088_ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__o211a_1
X_24118_ clknet_leaf_13_clk _00651_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24049_ clknet_leaf_34_clk _00582_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_16940_ _08870_ _09493_ _09495_ _09231_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__o211a_1
X_12063_ net559 _05045_ _05051_ _05049_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_1025 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16871_ _09211_ _09201_ VGND VGND VPWR VPWR _09428_ sky130_fd_sc_hd__and2_1
XFILLER_0_216_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18610_ _11033_ _11069_ VGND VGND VPWR VPWR _11070_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_205_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15822_ _08403_ _08402_ VGND VGND VPWR VPWR _08435_ sky130_fd_sc_hd__or2b_1
XFILLER_0_244_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19590_ _01374_ _01393_ _01420_ _01421_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__a211o_1
XTAP_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15753_ _08275_ _08315_ _08367_ VGND VGND VPWR VPWR _08368_ sky130_fd_sc_hd__o21ba_1
X_18541_ _10071_ _11001_ _11002_ _10620_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__o211a_1
X_12965_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _05759_ sky130_fd_sc_hd__clkbuf_4
XTAP_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14704_ _07390_ _07391_ _07342_ _07344_ VGND VGND VPWR VPWR _07393_ sky130_fd_sc_hd__o211ai_2
X_11916_ net717 _04964_ _04966_ _04955_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__o211a_1
XFILLER_0_185_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15684_ _08298_ _08299_ _08270_ _08271_ VGND VGND VPWR VPWR _08301_ sky130_fd_sc_hd__o211ai_1
X_18472_ _10587_ _10614_ _10612_ top_inst.grid_inst.data_path_wires\[12\]\[5\] VGND
+ VGND VPWR VPWR _10935_ sky130_fd_sc_hd__a22o_1
XTAP_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12896_ _05447_ _05306_ _05644_ _05700_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__o211a_1
XTAP_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _07319_ _07324_ VGND VGND VPWR VPWR _07325_ sky130_fd_sc_hd__xnor2_1
X_17423_ _09935_ _09956_ VGND VGND VPWR VPWR _09961_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_1091 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11847_ net282 _04925_ _04927_ _04916_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__o211a_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[24\] _09631_ VGND
+ VGND VPWR VPWR _09895_ sky130_fd_sc_hd__xnor2_1
X_14566_ net230 _07198_ _07256_ _07257_ VGND VGND VPWR VPWR _07258_ sky130_fd_sc_hd__a211oi_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11778_ top_inst.axis_out_inst.out_buff_data\[69\] _04877_ VGND VGND VPWR VPWR _04888_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_28_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_915 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16305_ _08677_ _08688_ _08884_ _08885_ VGND VGND VPWR VPWR _08887_ sky130_fd_sc_hd__nand4_4
X_13517_ _06265_ _06266_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__nand2_1
X_17285_ _08870_ _09828_ _09829_ _09231_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14497_ _05632_ _07190_ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_972 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16236_ _08794_ _08795_ _08818_ _08819_ VGND VGND VPWR VPWR _08820_ sky130_fd_sc_hd__a211oi_2
X_19024_ _11443_ _11444_ VGND VGND VPWR VPWR _11445_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13448_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _06208_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16167_ _08751_ _08752_ VGND VGND VPWR VPWR _08753_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13379_ _06120_ _06123_ _06151_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15118_ _07766_ _07764_ _07765_ VGND VGND VPWR VPWR _07768_ sky130_fd_sc_hd__and3_1
XFILLER_0_224_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16098_ _08669_ _08681_ _08691_ _08692_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19926_ _01720_ _01728_ _01744_ _01701_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__a22o_1
X_15049_ _07672_ _07679_ VGND VGND VPWR VPWR _07701_ sky130_fd_sc_hd__or2_1
XFILLER_0_220_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19857_ _01661_ _01663_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__nand2_1
XFILLER_0_236_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_235_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18808_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[3\]
+ top_inst.grid_inst.data_path_wires\[13\]\[2\] top_inst.grid_inst.data_path_wires\[13\]\[1\]
+ VGND VGND VPWR VPWR _11234_ sky130_fd_sc_hd__nand4_1
X_19788_ _01569_ _01581_ _01580_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_190_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18739_ net990 _10616_ _11169_ _11160_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_1347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21750_ _03278_ _03474_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20701_ _02477_ _02479_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21681_ _03407_ _03408_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_1130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23420_ _04869_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__buf_2
XFILLER_0_4_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20632_ _02363_ _02373_ _02412_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_163_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23351_ net512 _04791_ _04793_ _04782_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20563_ _02343_ _02345_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22302_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[18\]\[4\]
+ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23282_ net476 _04752_ _04754_ _04743_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__o211a_1
X_20494_ _01993_ _02229_ _02276_ _02277_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_1259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22233_ _03920_ _03921_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_203_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22164_ _03852_ _03853_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21115_ _02871_ _02869_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__or2_1
X_22095_ _03765_ _03768_ _03766_ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_61_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21046_ _02746_ _02786_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22997_ net971 _04588_ _04589_ _04590_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_241_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12750_ _05558_ _05559_ _05328_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__a21o_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21948_ _03662_ VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__clkbuf_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_733 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12681_ _05489_ _05491_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21879_ _03576_ _03597_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__xnor2_2
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _07116_ VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23618_ clknet_leaf_105_clk net574 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24598_ clknet_leaf_22_clk _01131_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_132_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_1327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14351_ net1042 _07048_ _07056_ _07058_ _06180_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__o221a_1
XFILLER_0_135_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23549_ clknet_leaf_131_clk _00082_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13302_ _06042_ _06038_ _06076_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__nand3_1
X_17070_ _09585_ _09614_ VGND VGND VPWR VPWR _09622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_181_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14282_ _06989_ _06992_ VGND VGND VPWR VPWR _06993_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_135_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16021_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[14\] _08452_ _08373_
+ VGND VGND VPWR VPWR _08629_ sky130_fd_sc_hd__a21o_1
X_13233_ top_inst.grid_inst.data_path_wires\[1\]\[4\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[6\]
+ _06008_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13164_ _05940_ _05942_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12115_ net469 _05071_ _05080_ _05075_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13095_ _05837_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__inv_2
X_17972_ _10473_ _10475_ VGND VGND VPWR VPWR _10476_ sky130_fd_sc_hd__xor2_1
X_19711_ _01537_ _01538_ _01532_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__a21oi_1
X_16923_ _09476_ _09477_ _09469_ VGND VGND VPWR VPWR _09479_ sky130_fd_sc_hd__a21o_1
X_12046_ net385 _05036_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19642_ _11722_ _01472_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__and2_1
X_16854_ _09367_ _09363_ VGND VGND VPWR VPWR _09411_ sky130_fd_sc_hd__or2b_1
XFILLER_0_233_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15805_ _08417_ _08418_ VGND VGND VPWR VPWR _08419_ sky130_fd_sc_hd__nor2_1
X_19573_ _11705_ _01403_ _01404_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__a21bo_1
X_16785_ _09331_ _09332_ _09342_ _09343_ VGND VGND VPWR VPWR _09344_ sky130_fd_sc_hd__nand4_2
X_13997_ _06628_ _06626_ _06640_ _06637_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__and4_1
XFILLER_0_232_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18524_ _10984_ _10985_ VGND VGND VPWR VPWR _10986_ sky130_fd_sc_hd__nand2_1
X_12948_ _05739_ _05567_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15736_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[7\] _08340_ VGND
+ VGND VPWR VPWR _08351_ sky130_fd_sc_hd__nand2_1
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18455_ _10917_ _10918_ VGND VGND VPWR VPWR _10919_ sky130_fd_sc_hd__and2_1
XFILLER_0_213_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12879_ _05658_ _05684_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__xnor2_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15667_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[5\] _08250_ _08251_
+ VGND VGND VPWR VPWR _08284_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17406_ _09933_ _09944_ VGND VGND VPWR VPWR _09945_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14618_ _07266_ _07268_ _07265_ VGND VGND VPWR VPWR _07309_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_28_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18386_ _10850_ VGND VGND VPWR VPWR _10851_ sky130_fd_sc_hd__inv_2
X_15598_ _08197_ _08217_ VGND VGND VPWR VPWR _08218_ sky130_fd_sc_hd__and2_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14549_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _07241_ sky130_fd_sc_hd__inv_2
X_17337_ _09872_ _09878_ VGND VGND VPWR VPWR _09879_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17268_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[19\] _09628_ _09629_
+ VGND VGND VPWR VPWR _09813_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19007_ _11413_ _11415_ VGND VGND VPWR VPWR _11428_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16219_ _08671_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[2\] _08800_
+ _08801_ VGND VGND VPWR VPWR _08803_ sky130_fd_sc_hd__nand4_2
XFILLER_0_114_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17199_ _08870_ _09746_ _09747_ _09231_ VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_1123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_220_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19909_ _01729_ _01730_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_209_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22920_ top_inst.skew_buff_inst.row\[2\].output_reg\[7\] _04543_ VGND VGND VPWR VPWR
+ _04546_ sky130_fd_sc_hd__or2_1
XFILLER_0_194_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22851_ net762 _04504_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21802_ _05405_ _03524_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__nor2_1
XFILLER_0_223_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22782_ _04449_ _04450_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_1263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24521_ clknet_leaf_128_clk _01054_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dfxtp_4
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21733_ _03420_ _03430_ _03454_ _03410_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_66_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24452_ clknet_leaf_64_clk _00985_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21664_ _03370_ _03391_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__or2_1
XFILLER_0_191_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23403_ net65 _04658_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20615_ _01999_ _02227_ _02368_ _02369_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__o2bb2ai_1
X_24383_ clknet_leaf_39_clk _00916_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21595_ _02895_ _03253_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23334_ net158 _04779_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20546_ _02003_ _02013_ _02011_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__and3_1
XFILLER_0_166_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_858 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23265_ net125 _04740_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__or2_1
X_20477_ _02260_ _02261_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22216_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[18\]\[2\]
+ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23196_ net92 _04701_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__or2_1
XTAP_6702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22147_ _03807_ _03808_ _03836_ _03837_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__a211o_1
XTAP_6724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22078_ _03739_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__inv_2
XTAP_6779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13920_ _05755_ VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__clkbuf_4
X_21029_ _02503_ _02785_ _02793_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__or3_1
XFILLER_0_195_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_215_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13851_ _06496_ _06591_ VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_241_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12802_ _05603_ _05608_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16570_ _09143_ _09144_ _08265_ VGND VGND VPWR VPWR _09146_ sky130_fd_sc_hd__o21a_1
X_13782_ _06196_ _06214_ _06524_ _06193_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_201_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12733_ _05494_ _05495_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__or2_1
X_15521_ _08152_ _08140_ VGND VGND VPWR VPWR _08153_ sky130_fd_sc_hd__or2_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15452_ _08092_ _08093_ VGND VGND VPWR VPWR _08094_ sky130_fd_sc_hd__nor2_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18240_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[5\] _09496_ _10707_
+ _10708_ VGND VGND VPWR VPWR _10709_ sky130_fd_sc_hd__a22o_1
X_12664_ _05441_ _05442_ _05474_ _05475_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__o211ai_4
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14403_ _07098_ _07099_ _07094_ VGND VGND VPWR VPWR _07101_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_203_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15383_ _08025_ _08026_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[12\]
+ _07816_ VGND VGND VPWR VPWR _08027_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_26_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18171_ _10626_ _10637_ VGND VGND VPWR VPWR _10642_ sky130_fd_sc_hd__or2b_1
X_12595_ _05376_ _05390_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17122_ _09213_ _09219_ _09597_ _09672_ VGND VGND VPWR VPWR _09673_ sky130_fd_sc_hd__a211o_1
X_14334_ _07041_ _07042_ VGND VGND VPWR VPWR _07043_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_243_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17053_ _09553_ _09561_ net1117 VGND VGND VPWR VPWR _09606_ sky130_fd_sc_hd__o21bai_1
X_14265_ _06974_ _06975_ VGND VGND VPWR VPWR _06976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_243_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_208_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16004_ _08570_ _08574_ _08572_ VGND VGND VPWR VPWR _08613_ sky130_fd_sc_hd__a21oi_2
X_13216_ _05943_ _05952_ _05993_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_243_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14196_ _06907_ _06908_ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13147_ top_inst.grid_inst.data_path_wires\[1\]\[1\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__and2b_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13078_ _05746_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[2\] _05857_
+ _05858_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__a22o_1
X_17955_ top_inst.grid_inst.data_path_wires\[11\]\[7\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _10459_ sky130_fd_sc_hd__nand2_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16906_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[9\] _09419_ VGND
+ VGND VPWR VPWR _09462_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12029_ _04911_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_174_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17886_ _10332_ _10348_ _10347_ VGND VGND VPWR VPWR _10392_ sky130_fd_sc_hd__o21bai_1
X_19625_ _01453_ _01454_ _01455_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__nand3_2
XFILLER_0_75_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16837_ _09346_ _09348_ VGND VGND VPWR VPWR _09395_ sky130_fd_sc_hd__and2b_1
XFILLER_0_220_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19556_ _01382_ _01383_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16768_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[6\] _09325_ _09326_
+ VGND VGND VPWR VPWR _09327_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18507_ _10968_ VGND VGND VPWR VPWR _10969_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15719_ _08333_ _08334_ VGND VGND VPWR VPWR _08335_ sky130_fd_sc_hd__xnor2_1
X_19487_ _01312_ _01319_ _01320_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__nand3_1
XFILLER_0_220_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16699_ _09259_ _09260_ VGND VGND VPWR VPWR _09261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18438_ _10900_ _10901_ VGND VGND VPWR VPWR _10902_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18369_ _10834_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20400_ top_inst.grid_inst.data_path_wires\[16\]\[7\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__nand2_2
XFILLER_0_173_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_1268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21380_ _03072_ _03112_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20331_ _01997_ _02007_ _02084_ _02083_ VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23050_ net5 _04615_ _04621_ _04619_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20262_ _01989_ _01986_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[3\]
+ _02051_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__nand4_1
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22001_ _03703_ _05275_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__or2_1
XTAP_6009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20193_ _10030_ _11696_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__or2_2
XFILLER_0_122_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23952_ clknet_leaf_90_clk _00485_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22903_ _02706_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__clkbuf_4
XTAP_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23883_ clknet_leaf_61_clk _00416_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22834_ _02706_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__buf_2
XFILLER_0_196_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_233_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22765_ _04426_ _04433_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24504_ clknet_leaf_128_clk _01037_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dfxtp_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21716_ top_inst.deskew_buff_inst.col_input\[82\] _03442_ _06140_ VGND VGND VPWR
+ VPWR _03443_ sky130_fd_sc_hd__mux2_1
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22696_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[23\] _04215_ _04216_
+ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_240_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24435_ clknet_leaf_54_clk _00968_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21647_ _03122_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__buf_4
XFILLER_0_30_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24366_ clknet_leaf_31_clk _00899_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[125\]
+ sky130_fd_sc_hd__dfxtp_1
X_12380_ net901 _05230_ _05231_ _05221_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_70 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21578_ net818 _02638_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__or2_1
XANTENNA_81 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_92 net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23317_ net150 _04766_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20529_ _02271_ _02302_ _02301_ VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_166_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24297_ clknet_leaf_137_clk _00830_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[72\]
+ sky130_fd_sc_hd__dfxtp_1
X_14050_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[6\] _05406_ VGND
+ VGND VPWR VPWR _06767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23248_ net117 _04727_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__or2_1
XFILLER_0_240_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13001_ _05784_ _05785_ _05336_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__o21ai_1
XTAP_6510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23179_ net84 _04687_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__or2_1
XTAP_6521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17740_ _10247_ _10248_ VGND VGND VPWR VPWR _10249_ sky130_fd_sc_hd__and2b_1
XTAP_6598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14952_ top_inst.grid_inst.data_path_wires\[6\]\[5\] VGND VGND VPWR VPWR _07619_
+ sky130_fd_sc_hd__buf_4
XFILLER_0_238_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13903_ top_inst.grid_inst.data_path_wires\[3\]\[7\] VGND VGND VPWR VPWR _06635_
+ sky130_fd_sc_hd__clkbuf_4
X_17671_ _10156_ _10157_ _10180_ _10181_ VGND VGND VPWR VPWR _10182_ sky130_fd_sc_hd__a211oi_2
X_14883_ _07535_ _07560_ _07565_ VGND VGND VPWR VPWR _07567_ sky130_fd_sc_hd__nor3_1
XFILLER_0_242_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19410_ _01236_ _01237_ _01244_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16622_ _09193_ VGND VGND VPWR VPWR _09194_ sky130_fd_sc_hd__clkbuf_4
X_13834_ _06544_ _06543_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19341_ top_inst.deskew_buff_inst.col_input\[2\] _11723_ _01178_ _01179_ VGND VGND
+ VPWR VPWR _01180_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16553_ _09055_ _09127_ VGND VGND VPWR VPWR _09129_ sky130_fd_sc_hd__and2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13765_ _06507_ _06508_ VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15504_ _08139_ _08140_ VGND VGND VPWR VPWR _08141_ sky130_fd_sc_hd__or2_1
X_12716_ _05505_ _05514_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__nand2_1
X_19272_ top_inst.skew_buff_inst.row\[3\].output_reg\[0\] top_inst.axis_in_inst.inbuf_bus\[24\]
+ net205 VGND VGND VPWR VPWR _11676_ sky130_fd_sc_hd__mux2_2
XFILLER_0_167_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16484_ _09019_ _09025_ _09018_ VGND VGND VPWR VPWR _09062_ sky130_fd_sc_hd__a21o_1
X_13696_ _06439_ _06441_ VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_214_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18223_ _10581_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[2\] _10672_
+ _10645_ _10608_ VGND VGND VPWR VPWR _10692_ sky130_fd_sc_hd__a32o_1
X_12647_ _05457_ _05458_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15435_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[13\] _07924_ _07844_
+ VGND VGND VPWR VPWR _08077_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15366_ _08004_ _08009_ VGND VGND VPWR VPWR _08010_ sky130_fd_sc_hd__xnor2_1
X_18154_ _10625_ _10626_ _06682_ VGND VGND VPWR VPWR _10627_ sky130_fd_sc_hd__a21o_1
X_12578_ _05357_ _05361_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17105_ _09653_ _09656_ VGND VGND VPWR VPWR _09657_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14317_ _06980_ _07010_ _07025_ VGND VGND VPWR VPWR _07026_ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15297_ _07820_ _07864_ _07904_ _07942_ VGND VGND VPWR VPWR _07943_ sky130_fd_sc_hd__a31o_1
X_18085_ net859 _10563_ _10576_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold307 top_inst.axis_out_inst.out_buff_data\[71\] VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold318 _00006_ VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__dlygate4sd3_1
X_17036_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[11\] _09419_ VGND
+ VGND VPWR VPWR _09589_ sky130_fd_sc_hd__nand2_1
X_14248_ _06848_ _06958_ _06959_ _06684_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__o211a_1
Xhold329 _00157_ VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14179_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[3\]\[4\]
+ _06890_ VGND VGND VPWR VPWR _06892_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ _11401_ _11408_ VGND VGND VPWR VPWR _11409_ sky130_fd_sc_hd__xor2_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _10404_ _10442_ VGND VGND VPWR VPWR _10443_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17869_ _10052_ _10050_ _10040_ VGND VGND VPWR VPWR _10375_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_205_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19608_ _01437_ _01438_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20880_ _02528_ _02644_ _02650_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__nand3_1
XFILLER_0_75_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_230_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19539_ _01369_ _01370_ _01362_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22550_ _04193_ _04228_ _04229_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_75_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21501_ _09787_ _03232_ _03233_ _03234_ _09806_ VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__o311a_1
XFILLER_0_88_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22481_ _03937_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__buf_4
XFILLER_0_185_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24220_ clknet_leaf_19_clk _00753_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21432_ _03163_ _03166_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_920 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24151_ clknet_leaf_18_clk _00684_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21363_ _03097_ _03099_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_140_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23102_ net284 _10541_ _04649_ _04643_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20314_ _01990_ _02016_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[5\]
+ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__nand3_2
X_24082_ clknet_leaf_111_clk _00615_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold830 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[11\] VGND
+ VGND VPWR VPWR net1012 sky130_fd_sc_hd__dlygate4sd3_1
X_21294_ _03032_ VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold841 top_inst.axis_out_inst.out_buff_data\[63\] VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold852 top_inst.axis_in_inst.inbuf_bus\[27\] VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23033_ net29 _04601_ _04611_ _04606_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold863 top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[1\] VGND VGND
+ VPWR VPWR net1045 sky130_fd_sc_hd__dlygate4sd3_1
X_20245_ _02033_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__inv_2
Xhold874 top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[2\] VGND VGND
+ VPWR VPWR net1056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[15\] VGND VGND
+ VPWR VPWR net1067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold896 top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[0\] VGND VGND
+ VPWR VPWR net1078 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20176_ net490 _01202_ _01983_ _01985_ _01863_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__o221a_1
XTAP_5127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_239_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23935_ clknet_leaf_81_clk _00468_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23866_ clknet_leaf_78_clk _00399_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11880_ net411 _04938_ _04946_ _04942_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22817_ _04449_ _04469_ _04482_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_233_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23797_ clknet_leaf_70_clk _00330_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_196_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13550_ top_inst.grid_inst.data_path_wires\[2\]\[3\] _06186_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _06299_ sky130_fd_sc_hd__nand4_2
XFILLER_0_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22748_ _04417_ _04418_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_976 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12501_ net950 _05314_ _05319_ _05308_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13481_ _06219_ _06223_ _06232_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__o21a_1
XFILLER_0_180_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22679_ _04329_ _04332_ _04350_ _04312_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_81_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15220_ _06848_ _07865_ _07867_ _07643_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24418_ clknet_leaf_57_clk net644 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12432_ net304 _05256_ _05259_ _05261_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_834 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15151_ _07797_ _07798_ _07749_ _07751_ VGND VGND VPWR VPWR _07800_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24349_ clknet_leaf_23_clk _00882_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[108\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12363_ _05142_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_69_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14102_ _06632_ _06643_ _06815_ _06816_ VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_200_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15082_ _07700_ _07702_ VGND VGND VPWR VPWR _07733_ sky130_fd_sc_hd__or2b_1
X_12294_ _05142_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_239_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_240_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14033_ _06624_ _06692_ _06712_ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__a21o_1
X_18910_ _11333_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_238_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19890_ top_inst.deskew_buff_inst.col_input\[18\] _01712_ _06140_ VGND VGND VPWR
+ VPWR _01713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18841_ top_inst.grid_inst.data_path_wires\[13\]\[6\] top_inst.grid_inst.data_path_wires\[13\]\[5\]
+ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _11266_ sky130_fd_sc_hd__nand4_1
XTAP_6340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18772_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[2\] _11179_ _11180_
+ VGND VGND VPWR VPWR _11200_ sky130_fd_sc_hd__a21boi_4
XTAP_6395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15984_ _08557_ _08525_ _08567_ VGND VGND VPWR VPWR _08593_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_234_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17723_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[7\] _10198_ _10199_
+ VGND VGND VPWR VPWR _10232_ sky130_fd_sc_hd__a21boi_2
XTAP_5683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14935_ _05736_ _07061_ VGND VGND VPWR VPWR _07607_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17654_ _10160_ _10164_ VGND VGND VPWR VPWR _10165_ sky130_fd_sc_hd__xor2_1
X_14866_ _07484_ _07483_ _07516_ VGND VGND VPWR VPWR _07551_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_216_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16605_ _09175_ _09178_ VGND VGND VPWR VPWR _09179_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_212_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13817_ _06196_ _06524_ _06557_ VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__nor3_1
X_17585_ _10086_ _10079_ _10098_ VGND VGND VPWR VPWR _10099_ sky130_fd_sc_hd__a21o_1
XFILLER_0_225_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14797_ _07445_ _07478_ VGND VGND VPWR VPWR _07483_ sky130_fd_sc_hd__or2b_4
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19324_ _11717_ _11718_ _11712_ VGND VGND VPWR VPWR _11719_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_57_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16536_ _09072_ _09074_ _09112_ VGND VGND VPWR VPWR _09113_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_128_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13748_ _06490_ _06491_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19255_ _11667_ _11668_ VGND VGND VPWR VPWR _11669_ sky130_fd_sc_hd__xnor2_1
X_16467_ _09040_ _09044_ VGND VGND VPWR VPWR _09045_ sky130_fd_sc_hd__xor2_1
X_13679_ _06377_ _06378_ _06374_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__or3b_1
XFILLER_0_186_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18206_ _10647_ _10654_ VGND VGND VPWR VPWR _10676_ sky130_fd_sc_hd__or2_1
X_15418_ _08019_ _08060_ VGND VGND VPWR VPWR _08061_ sky130_fd_sc_hd__xor2_2
XFILLER_0_13_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19186_ _11563_ _11566_ _11602_ VGND VGND VPWR VPWR _11603_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16398_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[10\] _08897_ VGND
+ VGND VPWR VPWR _08978_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18137_ _10612_ _10057_ VGND VGND VPWR VPWR _10613_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15349_ _07621_ _07640_ _07991_ VGND VGND VPWR VPWR _07993_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold104 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[24\] VGND
+ VGND VPWR VPWR net286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold115 _00929_ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18068_ _10547_ _10551_ VGND VGND VPWR VPWR _10568_ sky130_fd_sc_hd__nand2_1
Xhold126 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[28\] VGND
+ VGND VPWR VPWR net308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[17\] VGND
+ VGND VPWR VPWR net319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_956 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold148 _00282_ VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17019_ _09571_ _09572_ VGND VGND VPWR VPWR _09573_ sky130_fd_sc_hd__nor2_2
XFILLER_0_22_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold159 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[18\] VGND
+ VGND VPWR VPWR net341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20030_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[25\] _01764_ VGND
+ VGND VPWR VPWR _01846_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21981_ _02871_ _02877_ _03689_ _03660_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23720_ clknet_leaf_121_clk _00253_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_20932_ _02700_ _02701_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__xnor2_1
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_234_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23651_ clknet_leaf_122_clk _00184_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_230_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20863_ _02541_ _02570_ _02633_ _02635_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__o31a_1
XFILLER_0_166_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_234_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22602_ _04251_ _04260_ _04278_ _06734_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23582_ clknet_leaf_106_clk _00115_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20794_ _02532_ _02546_ _02564_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22533_ net508 _06169_ _04213_ _03929_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22464_ _04145_ _04146_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24203_ clknet_leaf_16_clk _00736_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21415_ _03083_ _03100_ _03150_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22395_ _04020_ _04021_ _04037_ _04036_ _04034_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__o32a_1
XFILLER_0_115_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24134_ clknet_leaf_0_clk _00667_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_21346_ _03075_ _03082_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24065_ clknet_leaf_83_clk _00598_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_60_1110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold660 top_inst.axis_out_inst.out_buff_data\[121\] VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__dlygate4sd3_1
X_21277_ _03010_ _03015_ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__xnor2_1
Xhold671 _00926_ VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__dlygate4sd3_1
X_23016_ _04600_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__buf_4
Xhold682 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[18\] VGND
+ VGND VPWR VPWR net864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[11\] VGND
+ VGND VPWR VPWR net875 sky130_fd_sc_hd__dlygate4sd3_1
X_20228_ _02001_ _11163_ _02022_ _02006_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_217_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20159_ _01966_ _01968_ _10831_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__o21a_1
XTAP_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _05770_ sky130_fd_sc_hd__buf_2
XTAP_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14720_ _07406_ _07407_ VGND VGND VPWR VPWR _07408_ sky130_fd_sc_hd__xnor2_1
XTAP_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23918_ clknet_leaf_77_clk _00451_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ net880 _04964_ _04975_ _04968_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__o211a_1
XTAP_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14651_ _07332_ _07340_ VGND VGND VPWR VPWR _07341_ sky130_fd_sc_hd__xor2_1
XTAP_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ net924 _04925_ _04936_ _04929_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23849_ clknet_leaf_95_clk _00382_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _06340_ _06349_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__xor2_1
XFILLER_0_200_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17370_ _09902_ _09903_ VGND VGND VPWR VPWR _09910_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ _07232_ _07228_ VGND VGND VPWR VPWR _07273_ sky130_fd_sc_hd__or2b_1
XFILLER_0_170_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11794_ net705 _04890_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16321_ _08893_ _08849_ _08901_ VGND VGND VPWR VPWR _08903_ sky130_fd_sc_hd__nor3_1
XFILLER_0_27_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13533_ _06235_ _06257_ _06282_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19040_ _11420_ _11459_ VGND VGND VPWR VPWR _11461_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16252_ _08833_ _08834_ VGND VGND VPWR VPWR _08835_ sky130_fd_sc_hd__xnor2_1
X_13464_ net1017 _05788_ _06218_ _06207_ VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_207_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15203_ _07841_ _07797_ _07849_ VGND VGND VPWR VPWR _07851_ sky130_fd_sc_hd__nor3_1
X_12415_ net333 _05243_ _05251_ _05247_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16183_ _08669_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[2\] VGND
+ VGND VPWR VPWR _08768_ sky130_fd_sc_hd__nand2_1
X_13395_ _06167_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15134_ _07781_ _07782_ VGND VGND VPWR VPWR _07783_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12346_ net698 _05204_ _05212_ _05208_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19942_ _01396_ VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__clkbuf_4
X_15065_ _07714_ _07715_ VGND VGND VPWR VPWR _07716_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12277_ net306 _05169_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14016_ _06733_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19873_ net1096 _01202_ _01695_ _01696_ _11228_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__o221a_1
XFILLER_0_219_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18824_ _11247_ _11249_ VGND VGND VPWR VPWR _11250_ sky130_fd_sc_hd__xnor2_2
XTAP_6170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_234_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18755_ _11182_ _11183_ VGND VGND VPWR VPWR _11184_ sky130_fd_sc_hd__xnor2_1
XTAP_5480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15967_ _08568_ _08569_ _08575_ VGND VGND VPWR VPWR _08577_ sky130_fd_sc_hd__a21oi_1
XTAP_5491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17706_ _10209_ _10215_ VGND VGND VPWR VPWR _10216_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14918_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[19\] _07595_ VGND
+ VGND VPWR VPWR _07598_ sky130_fd_sc_hd__and2_1
XFILLER_0_175_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18686_ top_inst.grid_inst.data_path_wires\[13\]\[1\] VGND VGND VPWR VPWR _11132_
+ sky130_fd_sc_hd__clkbuf_4
XTAP_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15898_ _08478_ _08479_ _08508_ VGND VGND VPWR VPWR _08510_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17637_ _10146_ _10148_ VGND VGND VPWR VPWR _10149_ sky130_fd_sc_hd__xor2_1
X_14849_ _07532_ _07533_ VGND VGND VPWR VPWR _07534_ sky130_fd_sc_hd__or2b_1
XFILLER_0_188_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17568_ net1036 VGND VGND VPWR VPWR _10083_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19307_ _11704_ VGND VGND VPWR VPWR _11705_ sky130_fd_sc_hd__buf_2
XFILLER_0_163_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16519_ _09055_ _09094_ VGND VGND VPWR VPWR _09096_ sky130_fd_sc_hd__and2_1
XFILLER_0_175_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17499_ top_inst.grid_inst.data_path_wires\[11\]\[3\] VGND VGND VPWR VPWR _10029_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19238_ _11624_ _11627_ _11652_ VGND VGND VPWR VPWR _11653_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_186_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19169_ _11551_ _11555_ _11553_ VGND VGND VPWR VPWR _11586_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21200_ _05312_ _02939_ _02940_ _02941_ VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22180_ _03866_ _03869_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_223_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21131_ _02883_ _02021_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1098 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21062_ _02807_ _02809_ _02826_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_111_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20013_ _01561_ _01829_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__xor2_2
XFILLER_0_226_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_216_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21964_ _03663_ _03664_ _03671_ _03676_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20915_ _02656_ _02680_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__nor2_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23703_ clknet_leaf_116_clk _00236_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21895_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[27\] _03376_ VGND
+ VGND VPWR VPWR _03613_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23634_ clknet_leaf_125_clk net931 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20846_ _02466_ _02617_ _02618_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23565_ clknet_leaf_100_clk net721 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20777_ _02551_ _02552_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22516_ _04061_ _04195_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23496_ clknet_leaf_140_clk net475 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[86\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22447_ _04061_ _04128_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12200_ _05009_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__buf_2
XFILLER_0_66_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13180_ _05956_ _05958_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__xnor2_1
X_22378_ _04061_ _04062_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12131_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[28\] _05089_
+ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__or2_1
X_24117_ clknet_leaf_12_clk _00650_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_21329_ _03064_ _03065_ _05353_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24048_ clknet_leaf_34_clk _00581_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12062_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[30\] _05050_
+ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__or2_1
Xhold490 top_inst.deskew_buff_inst.col_input\[54\] VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16870_ _09423_ _09426_ VGND VGND VPWR VPWR _09427_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15821_ net1086 _07048_ _08433_ _08434_ _07708_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__o221a_1
XFILLER_0_244_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_232_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18540_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[12\] _10639_ VGND
+ VGND VPWR VPWR _11002_ sky130_fd_sc_hd__or2_1
XFILLER_0_232_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15752_ _08316_ _08319_ _08320_ VGND VGND VPWR VPWR _08367_ sky130_fd_sc_hd__and3_1
XTAP_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _05734_ _05756_ _05758_ _05743_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__o211a_1
XTAP_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14703_ _07342_ _07344_ _07390_ _07391_ VGND VGND VPWR VPWR _07392_ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11915_ net493 _04956_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__or2_1
XTAP_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18471_ _10589_ _10587_ _10614_ _10612_ VGND VGND VPWR VPWR _10934_ sky130_fd_sc_hd__and4_1
XFILLER_0_217_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _08270_ _08271_ _08298_ _08299_ VGND VGND VPWR VPWR _08300_ sky130_fd_sc_hd__a211o_1
XTAP_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _05302_ _05306_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__nand2_1
XTAP_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _09958_ _09959_ VGND VGND VPWR VPWR _09960_ sky130_fd_sc_hd__nor2_1
X_14634_ _07322_ _07323_ VGND VGND VPWR VPWR _07324_ sky130_fd_sc_hd__nor2_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11846_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[2\] _04917_
+ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__or2_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17353_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[23\] _09628_ _09629_
+ VGND VGND VPWR VPWR _09894_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ _07253_ _07254_ _07255_ VGND VGND VPWR VPWR _07257_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11777_ net348 _04885_ _04887_ _04875_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _08677_ _08688_ _08884_ _08885_ VGND VGND VPWR VPWR _08886_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13516_ top_inst.grid_inst.data_path_wires\[2\]\[2\] _06184_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _06266_ sky130_fd_sc_hd__nand4_1
X_17284_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[20\] _09494_ VGND
+ VGND VPWR VPWR _09829_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_927 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14496_ _07160_ _07189_ _05316_ VGND VGND VPWR VPWR _07190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19023_ _11164_ top_inst.grid_inst.data_path_wires\[13\]\[4\] top_inst.grid_inst.data_path_wires\[13\]\[3\]
+ _11351_ VGND VGND VPWR VPWR _11444_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_36_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16235_ _08817_ _08815_ _08816_ VGND VGND VPWR VPWR _08819_ sky130_fd_sc_hd__and3_1
XFILLER_0_181_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13447_ _06186_ _06204_ _06206_ _06207_ VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16166_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[8\]\[1\]
+ top_inst.grid_inst.data_path_wires\[8\]\[0\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[4\]
+ VGND VGND VPWR VPWR _08752_ sky130_fd_sc_hd__a22o_1
X_13378_ _06054_ _06150_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15117_ _07764_ _07765_ _07766_ VGND VGND VPWR VPWR _07767_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12329_ net586 _05191_ _05202_ _05195_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__o211a_1
XFILLER_0_220_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16097_ _07617_ VGND VGND VPWR VPWR _08692_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_224_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19925_ _01737_ _01745_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__xnor2_1
X_15048_ _07695_ _07699_ VGND VGND VPWR VPWR _07700_ sky130_fd_sc_hd__xor2_2
XFILLER_0_103_1025 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19856_ _01668_ _01656_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18807_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[13\]\[2\]
+ top_inst.grid_inst.data_path_wires\[13\]\[1\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[4\]
+ VGND VGND VPWR VPWR _11233_ sky130_fd_sc_hd__a22o_1
XFILLER_0_235_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19787_ _01603_ _01613_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__xnor2_1
X_16999_ _09551_ _09552_ VGND VGND VPWR VPWR _09553_ sky130_fd_sc_hd__nand2_2
XFILLER_0_155_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18738_ _11167_ _11168_ _08181_ VGND VGND VPWR VPWR _11169_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_91_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18669_ _11117_ _11125_ VGND VGND VPWR VPWR _11126_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_222_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20700_ _02436_ _02442_ _02478_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__a21o_1
XFILLER_0_231_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21680_ _03246_ _03406_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__and2_1
XFILLER_0_188_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20631_ _02372_ _02371_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__and2b_1
XFILLER_0_50_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23350_ net39 _04792_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__or2_1
X_20562_ _02264_ _02308_ _02344_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_73_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22301_ top_inst.grid_inst.data_path_wires\[18\]\[3\] top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__and2b_1
X_23281_ net133 _04753_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__or2_1
X_20493_ top_inst.grid_inst.data_path_wires\[16\]\[5\] _02015_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[9\]
+ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__and3_1
XFILLER_0_144_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22232_ _03875_ _03848_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__or2b_1
XFILLER_0_30_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22163_ _03695_ _03693_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[1\]
+ _03697_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__nand4_1
XFILLER_0_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21114_ top_inst.grid_inst.data_path_wires\[17\]\[4\] VGND VGND VPWR VPWR _02871_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_1351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22094_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[4\] _03758_ _03759_
+ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_121_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21045_ _02799_ _02798_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__or2b_1
XFILLER_0_201_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22996_ _04550_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__buf_4
XFILLER_0_213_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21947_ _03311_ _03661_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__and2_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _05447_ _05449_ _05279_ _05490_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__or4_1
XFILLER_0_167_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21878_ _03596_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__inv_2
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23617_ clknet_leaf_105_clk net588 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_20829_ _02517_ _02595_ _02602_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24597_ clknet_leaf_22_clk _01130_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_126_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14350_ _07050_ _07055_ _07057_ VGND VGND VPWR VPWR _07058_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23548_ clknet_leaf_130_clk _00081_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13301_ _06042_ _06038_ _06076_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14281_ _06990_ _06957_ _06991_ VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23479_ clknet_leaf_134_clk net363 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13232_ _05746_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[6\] _06008_
+ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__a21oi_1
X_16020_ _08484_ _08598_ VGND VGND VPWR VPWR _08628_ sky130_fd_sc_hd__and2b_1
XFILLER_0_165_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13163_ _05855_ _05893_ _05941_ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_62_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12114_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[21\] _05076_
+ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__or2_1
XFILLER_0_237_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13094_ _05849_ _05850_ _05873_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__and3_1
X_17971_ _10418_ _10433_ _10474_ VGND VGND VPWR VPWR _10475_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19710_ _01532_ _01537_ _01538_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__and3_1
X_16922_ _09469_ _09476_ _09477_ VGND VGND VPWR VPWR _09478_ sky130_fd_sc_hd__nand3_1
X_12045_ net647 _05031_ _05040_ _05035_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19641_ top_inst.deskew_buff_inst.col_input\[10\] _11723_ _01470_ _01471_ VGND VGND
+ VPWR VPWR _01472_ sky130_fd_sc_hd__a22o_1
XFILLER_0_217_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16853_ _09391_ _09393_ VGND VGND VPWR VPWR _09410_ sky130_fd_sc_hd__nor2_2
XFILLER_0_233_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15804_ _08362_ _08364_ _08416_ VGND VGND VPWR VPWR _08418_ sky130_fd_sc_hd__and3_1
X_19572_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[4\] net195 _11704_
+ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _01404_ sky130_fd_sc_hd__a22o_1
XFILLER_0_233_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16784_ _09340_ _09341_ _09308_ VGND VGND VPWR VPWR _09343_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13996_ _06708_ _06713_ VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_87_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18523_ _10933_ _10983_ VGND VGND VPWR VPWR _10985_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15735_ _08339_ _08338_ VGND VGND VPWR VPWR _08350_ sky130_fd_sc_hd__or2b_1
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12947_ top_inst.grid_inst.data_path_wires\[1\]\[4\] VGND VGND VPWR VPWR _05746_
+ sky130_fd_sc_hd__clkbuf_4
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_1430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ _10881_ _10916_ VGND VGND VPWR VPWR _10918_ sky130_fd_sc_hd__or2_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15666_ _08245_ _08282_ VGND VGND VPWR VPWR _08283_ sky130_fd_sc_hd__xor2_1
X_12878_ _05682_ _05683_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__xor2_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17405_ _09942_ _09943_ VGND VGND VPWR VPWR _09944_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ _07306_ _07307_ VGND VGND VPWR VPWR _07308_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18385_ top_inst.grid_inst.data_path_wires\[12\]\[6\] top_inst.grid_inst.data_path_wires\[12\]\[5\]
+ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _10850_ sky130_fd_sc_hd__and4_1
X_11829_ net694 _04917_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__or2_1
XFILLER_0_233_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15597_ _05887_ _08214_ _08215_ _08216_ VGND VGND VPWR VPWR _08217_ sky130_fd_sc_hd__a31o_1
XFILLER_0_145_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17336_ _09877_ _09869_ VGND VGND VPWR VPWR _09878_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_776 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14548_ _07236_ _07239_ VGND VGND VPWR VPWR _07240_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17267_ _09792_ _09794_ _09811_ VGND VGND VPWR VPWR _09812_ sky130_fd_sc_hd__a21o_1
X_14479_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[2\] _07073_ _07171_
+ _07172_ VGND VGND VPWR VPWR _07173_ sky130_fd_sc_hd__nand4_2
XFILLER_0_148_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19006_ _11383_ _11422_ _11426_ _11382_ VGND VGND VPWR VPWR _11427_ sky130_fd_sc_hd__a22o_1
XFILLER_0_226_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16218_ _08671_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[2\] _08800_
+ _08801_ VGND VGND VPWR VPWR _08802_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17198_ net1080 _09494_ VGND VGND VPWR VPWR _09747_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16149_ _08723_ _08717_ _08735_ VGND VGND VPWR VPWR _08736_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_1135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19908_ _01697_ _01703_ _01727_ _01688_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_209_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19839_ _01661_ _01662_ _01658_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__a21o_1
XFILLER_0_236_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22850_ net987 _04496_ _04506_ _04498_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21801_ _03522_ _03523_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22781_ _04192_ _04431_ _04448_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24520_ clknet_leaf_132_clk _01053_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dfxtp_4
X_21732_ _03456_ _03457_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24451_ clknet_leaf_63_clk _00984_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21663_ _03370_ _03391_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23402_ net410 _04655_ _04821_ _04819_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__o211a_1
X_20614_ _02358_ _02360_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__or2_1
X_24382_ clknet_leaf_38_clk _00915_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21594_ _03253_ _03323_ _03324_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23333_ net434 _04778_ _04783_ _04782_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__o211a_1
X_20545_ _02013_ _02011_ _02003_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_140_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_140_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_127_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1008 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23264_ net730 _04739_ _04744_ _04743_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20476_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[7\] _02211_ _02210_
+ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_160_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22215_ top_inst.grid_inst.data_path_wires\[18\]\[1\] _03713_ VGND VGND VPWR VPWR
+ _03904_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23195_ net493 _04700_ _04705_ _04704_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22146_ _03834_ _03835_ _03809_ _03810_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__o211a_1
XTAP_6714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22077_ _03764_ _03769_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__xnor2_2
XTAP_6769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21028_ _02503_ _02785_ _02793_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_22_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13850_ _06588_ _06589_ _06590_ VGND VGND VPWR VPWR _06591_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_88_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12801_ _05603_ _05608_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__or2_1
XFILLER_0_241_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13781_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _06524_ sky130_fd_sc_hd__inv_2
X_22979_ top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[0\] _04570_ VGND
+ VGND VPWR VPWR _04580_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15520_ top_inst.grid_inst.data_path_wires\[7\]\[7\] VGND VGND VPWR VPWR _08152_
+ sky130_fd_sc_hd__buf_4
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12732_ _05540_ _05541_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__nand2_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_214_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_721 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15451_ _08058_ _08091_ VGND VGND VPWR VPWR _08093_ sky130_fd_sc_hd__and2_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12663_ _05472_ _05473_ _05443_ _05429_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__a211o_1
XFILLER_0_155_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14402_ _07098_ _07099_ _07094_ VGND VGND VPWR VPWR _07100_ sky130_fd_sc_hd__o21ba_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18170_ _04873_ VGND VGND VPWR VPWR _10641_ sky130_fd_sc_hd__buf_2
XFILLER_0_154_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15382_ _08022_ _08024_ _06404_ VGND VGND VPWR VPWR _08026_ sky130_fd_sc_hd__a21o_1
X_12594_ _05394_ _05396_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17121_ _09361_ _09219_ VGND VGND VPWR VPWR _09672_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14333_ _07039_ _07040_ VGND VGND VPWR VPWR _07042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_131_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_131_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_145_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17052_ _09602_ _09603_ _09553_ VGND VGND VPWR VPWR _09605_ sky130_fd_sc_hd__o21ai_1
X_14264_ _06961_ _06962_ _06973_ VGND VGND VPWR VPWR _06975_ sky130_fd_sc_hd__nand3_1
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16003_ _08610_ _08611_ VGND VGND VPWR VPWR _08612_ sky130_fd_sc_hd__nand2_1
X_13215_ _05942_ _05940_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__and2b_1
XFILLER_0_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14195_ _06825_ _06906_ VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13146_ _05918_ _05916_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ top_inst.grid_inst.data_path_wires\[1\]\[3\] _05741_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _05858_ sky130_fd_sc_hd__nand4_2
X_17954_ _10423_ _10424_ _10426_ VGND VGND VPWR VPWR _10458_ sky130_fd_sc_hd__or3_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16905_ _09198_ _09215_ _09426_ _09425_ VGND VGND VPWR VPWR _09461_ sky130_fd_sc_hd__a31o_1
X_12028_ net270 _05018_ _05030_ _05022_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17885_ _10374_ _10390_ VGND VGND VPWR VPWR _10391_ sky130_fd_sc_hd__xor2_1
XFILLER_0_178_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_217_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16836_ _09391_ _09392_ _09329_ _09331_ VGND VGND VPWR VPWR _09394_ sky130_fd_sc_hd__o211a_1
X_19624_ _01406_ _01414_ _01413_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_232_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_233_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19555_ _11177_ _01385_ _01387_ _11714_ VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__o211a_1
X_16767_ _09193_ _09188_ _09210_ net202 VGND VGND VPWR VPWR _09326_ sky130_fd_sc_hd__nand4_1
XFILLER_0_177_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13979_ _06675_ _06697_ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__xnor2_1
X_18506_ _10853_ _10931_ _10892_ VGND VGND VPWR VPWR _10968_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_244_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_244_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15718_ _08245_ _08282_ _08293_ VGND VGND VPWR VPWR _08334_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_244_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19486_ _01317_ _01318_ _01275_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__a21o_1
X_16698_ _09247_ _09240_ _09257_ VGND VGND VPWR VPWR _09260_ sky130_fd_sc_hd__or3_1
XFILLER_0_158_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18437_ _10855_ _10858_ _10856_ VGND VGND VPWR VPWR _10901_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_185_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15649_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[5\] _08066_ _08264_
+ _08266_ VGND VGND VPWR VPWR _08267_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18368_ _10641_ _10833_ VGND VGND VPWR VPWR _10834_ sky130_fd_sc_hd__and2_1
XFILLER_0_173_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17319_ _09844_ _09860_ VGND VGND VPWR VPWR _09862_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18299_ _10764_ _10765_ VGND VGND VPWR VPWR _10766_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_122_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20330_ _02115_ _02116_ _02108_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_998 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20261_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _02051_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22000_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _03703_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20192_ top_inst.grid_inst.data_path_wires\[16\]\[4\] VGND VGND VPWR VPWR _01997_
+ sky130_fd_sc_hd__buf_4
XFILLER_0_196_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_719 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23951_ clknet_leaf_90_clk _00484_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22902_ top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[7\] _04530_ VGND
+ VGND VPWR VPWR _04536_ sky130_fd_sc_hd__or2_1
XTAP_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23882_ clknet_leaf_63_clk _00415_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22833_ top_inst.skew_buff_inst.row\[3\].output_reg\[1\] _03691_ VGND VGND VPWR VPWR
+ _04497_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_224_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22764_ _04426_ _04433_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24503_ clknet_leaf_127_clk _01036_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21715_ _03438_ _03441_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22695_ _04343_ _04347_ _04346_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__a21o_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24434_ clknet_leaf_58_clk _00967_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_21646_ _03374_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__buf_2
XFILLER_0_168_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_951 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24365_ clknet_leaf_31_clk _00898_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[124\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21577_ _03277_ _03308_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_113_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_60 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_71 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_82 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23316_ net391 _04765_ _04773_ _04769_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__o211a_1
X_20528_ _02305_ _02306_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24296_ clknet_leaf_137_clk _00829_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23247_ net945 _04726_ _04734_ _04730_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__o211a_1
X_20459_ _02241_ _02242_ _02243_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13000_ _05734_ _05761_ _05783_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23178_ net548 _04685_ _04695_ _04691_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__o211a_1
XTAP_6511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22129_ _03812_ _03819_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__xnor2_1
XTAP_6544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14951_ _07615_ _07611_ _07616_ _07618_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__o211a_1
XTAP_6599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13902_ _05177_ VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__clkbuf_4
XTAP_5887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17670_ _10178_ _10179_ _10158_ VGND VGND VPWR VPWR _10181_ sky130_fd_sc_hd__a21oi_1
X_14882_ _07535_ _07560_ _07565_ VGND VGND VPWR VPWR _07566_ sky130_fd_sc_hd__o21a_1
XTAP_5898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16621_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _09193_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_173_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13833_ _06555_ _06574_ VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_203_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_230_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19340_ net172 _11732_ _10831_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16552_ _09055_ _09127_ VGND VGND VPWR VPWR _09128_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13764_ _06385_ _06506_ VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__and2_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_1123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15503_ _06619_ VGND VGND VPWR VPWR _08140_ sky130_fd_sc_hd__buf_2
XFILLER_0_210_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12715_ _05502_ _05504_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__or2_1
X_19271_ net748 _11662_ _11675_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16483_ _09053_ _09060_ VGND VGND VPWR VPWR _09061_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13695_ _06396_ _06398_ _06440_ VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__o21a_1
XFILLER_0_210_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18222_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[4\] _10664_ _10665_
+ VGND VGND VPWR VPWR _10691_ sky130_fd_sc_hd__a21boi_2
X_15434_ _08074_ _08075_ VGND VGND VPWR VPWR _08076_ sky130_fd_sc_hd__or2b_1
X_12646_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[2\] _05297_ VGND
+ VGND VPWR VPWR _05458_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18153_ _10617_ _10623_ _10624_ VGND VGND VPWR VPWR _10626_ sky130_fd_sc_hd__nand3_2
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15365_ _08007_ _08008_ VGND VGND VPWR VPWR _08009_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_104_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12577_ _05376_ _05390_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__xor2_1
XFILLER_0_182_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17104_ _09654_ _09655_ VGND VGND VPWR VPWR _09656_ sky130_fd_sc_hd__nand2_1
X_14316_ _07007_ _07009_ VGND VGND VPWR VPWR _07025_ sky130_fd_sc_hd__or2b_1
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18084_ net1076 _10563_ _10576_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__o21a_1
XFILLER_0_230_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15296_ _07869_ _07862_ _07903_ VGND VGND VPWR VPWR _07942_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold308 top_inst.deskew_buff_inst.col_input\[31\] VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17035_ _09194_ _09189_ _09219_ VGND VGND VPWR VPWR _09588_ sky130_fd_sc_hd__nand3_2
XFILLER_0_145_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold319 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[17\] VGND
+ VGND VPWR VPWR net501 sky130_fd_sc_hd__dlygate4sd3_1
X_14247_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[11\] _06168_ VGND
+ VGND VPWR VPWR _06959_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14178_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[6\] _06628_ _06890_
+ VGND VGND VPWR VPWR _06891_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13129_ _05902_ _05908_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__xnor2_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18986_ _11406_ _11407_ VGND VGND VPWR VPWR _11408_ sky130_fd_sc_hd__xnor2_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17937_ _10397_ _10441_ VGND VGND VPWR VPWR _10442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1035 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17868_ _10368_ _10373_ VGND VGND VPWR VPWR _10374_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_205_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19607_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[10\] _01354_ VGND
+ VGND VPWR VPWR _01438_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16819_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _09377_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17799_ _10290_ _10291_ _10306_ VGND VGND VPWR VPWR _10307_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_220_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19538_ _01362_ _01369_ _01370_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__nand3_1
XFILLER_0_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19469_ _11684_ _01301_ _01302_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21500_ net753 _05316_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22480_ _04137_ _04141_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21431_ _03164_ _03165_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_146_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24150_ clknet_leaf_18_clk _00683_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21362_ _03049_ _03055_ _03098_ VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__o21a_1
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23101_ top_inst.valid_pipe\[4\] _05323_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20313_ _02089_ _02090_ _02088_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__or3b_1
XFILLER_0_86_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24081_ clknet_leaf_111_clk _00614_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold820 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[20\] VGND VGND
+ VPWR VPWR net1002 sky130_fd_sc_hd__dlygate4sd3_1
X_21293_ _02135_ _03031_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold831 top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[8\] VGND VGND
+ VPWR VPWR net1013 sky130_fd_sc_hd__dlygate4sd3_1
X_23032_ top_inst.axis_in_inst.inbuf_bus\[6\] _04603_ VGND VGND VPWR VPWR _04611_
+ sky130_fd_sc_hd__or2_1
Xhold842 top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[9\] VGND VGND
+ VPWR VPWR net1024 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold853 top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[15\] VGND VGND
+ VPWR VPWR net1035 sky130_fd_sc_hd__dlygate4sd3_1
X_20244_ net760 _01735_ _02034_ _02035_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold864 top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[21\] VGND VGND
+ VPWR VPWR net1046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[25\] VGND VGND
+ VPWR VPWR net1057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_228_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold886 top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[0\] VGND VGND
+ VPWR VPWR net1068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold897 top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[2\] VGND VGND
+ VPWR VPWR net1079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20175_ _01964_ _01969_ _01982_ _01984_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__a31o_1
XTAP_5106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23934_ clknet_leaf_81_clk _00467_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_1392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23865_ clknet_leaf_68_clk _00398_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22816_ _04445_ _04481_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_212_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23796_ clknet_leaf_69_clk _00329_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_233_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22747_ _04386_ _04397_ _04413_ _04374_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12500_ _05317_ _05318_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13480_ top_inst.grid_inst.data_path_wires\[2\]\[3\] top_inst.grid_inst.data_path_wires\[2\]\[2\]
+ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__and4_1
XFILLER_0_192_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22678_ _04344_ _04351_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24417_ clknet_leaf_56_clk _00950_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12431_ _05260_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__buf_6
XFILLER_0_125_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21629_ _03349_ _03350_ _03358_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15150_ _07749_ _07751_ _07797_ _07798_ VGND VGND VPWR VPWR _07799_ sky130_fd_sc_hd__a211oi_2
X_24348_ clknet_leaf_24_clk _00881_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[107\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12362_ net929 _05217_ _05220_ _05221_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14101_ top_inst.grid_inst.data_path_wires\[3\]\[5\] _06648_ _06628_ _06645_ VGND
+ VGND VPWR VPWR _06816_ sky130_fd_sc_hd__nand4_1
XFILLER_0_240_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15081_ _07729_ _07731_ VGND VGND VPWR VPWR _07732_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12293_ net642 _05178_ _05181_ _05182_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24279_ clknet_leaf_11_clk _00812_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[17\]\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_14032_ _06739_ _06748_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_240_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18840_ top_inst.grid_inst.data_path_wires\[13\]\[5\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[13\]\[6\]
+ VGND VGND VPWR VPWR _11265_ sky130_fd_sc_hd__a22o_1
XTAP_6330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18771_ _11197_ _11198_ VGND VGND VPWR VPWR _11199_ sky130_fd_sc_hd__or2_1
XTAP_5640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15983_ _08556_ _08592_ _05440_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__a21oi_1
XTAP_6385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17722_ _10196_ _10202_ _10230_ VGND VGND VPWR VPWR _10231_ sky130_fd_sc_hd__a21o_1
XTAP_5673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14934_ top_inst.grid_inst.data_path_wires\[6\]\[0\] VGND VGND VPWR VPWR _07606_
+ sky130_fd_sc_hd__clkbuf_4
XTAP_5684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[6\] _10163_ VGND
+ VGND VPWR VPWR _10164_ sky130_fd_sc_hd__xor2_2
XFILLER_0_76_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14865_ _07548_ _07549_ VGND VGND VPWR VPWR _07550_ sky130_fd_sc_hd__and2_1
XFILLER_0_199_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16604_ _09163_ _09177_ VGND VGND VPWR VPWR _09178_ sky130_fd_sc_hd__xnor2_1
X_13816_ _06196_ _06524_ _06557_ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__o21a_1
X_17584_ _10090_ _10097_ VGND VGND VPWR VPWR _10098_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14796_ net1065 _06660_ _07482_ _07092_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19323_ _11715_ _11716_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[1\]
+ VGND VGND VPWR VPWR _11718_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16535_ _09032_ _09071_ VGND VGND VPWR VPWR _09112_ sky130_fd_sc_hd__and2b_1
XFILLER_0_161_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13747_ _06451_ _06454_ _06452_ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_168_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19254_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[16\] _11387_ _11338_
+ VGND VGND VPWR VPWR _11668_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_183_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16466_ _09042_ _09043_ VGND VGND VPWR VPWR _09044_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13678_ _06373_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18205_ _10670_ _10674_ VGND VGND VPWR VPWR _10675_ sky130_fd_sc_hd__xor2_2
X_15417_ _08058_ _08059_ VGND VGND VPWR VPWR _08060_ sky130_fd_sc_hd__and2_1
X_12629_ _05411_ _05431_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19185_ _11479_ _11601_ VGND VGND VPWR VPWR _11602_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_241_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16397_ _08679_ _08688_ _08928_ _08929_ VGND VGND VPWR VPWR _08977_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_207_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18136_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _10612_ sky130_fd_sc_hd__buf_2
XFILLER_0_186_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15348_ _07621_ _07640_ _07991_ VGND VGND VPWR VPWR _07992_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18067_ _10413_ _10549_ _10566_ VGND VGND VPWR VPWR _10567_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold105 _00287_ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15279_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[9\] _07924_ _07844_
+ VGND VGND VPWR VPWR _07925_ sky130_fd_sc_hd__a21o_1
Xhold116 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[21\] VGND
+ VGND VPWR VPWR net298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold127 _00195_ VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold138 _00280_ VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ _09569_ _09570_ _09542_ VGND VGND VPWR VPWR _09572_ sky130_fd_sc_hd__a21oi_1
Xhold149 top_inst.valid_pipe\[6\] VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18969_ _11345_ _11347_ _11389_ VGND VGND VPWR VPWR _11391_ sky130_fd_sc_hd__and3_1
XFILLER_0_226_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21980_ _03688_ _02869_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__or2_1
XFILLER_0_241_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20931_ _02673_ _02676_ _02671_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__o21a_1
XFILLER_0_221_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23650_ clknet_leaf_132_clk net347 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_20862_ _02569_ _02633_ _02634_ _02610_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_1140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22601_ _04251_ _04260_ _04278_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_194_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23581_ clknet_leaf_107_clk _00114_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_20793_ net268 _05634_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22532_ _04211_ _04212_ _05732_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22463_ _04097_ _04098_ _04111_ _04110_ _04108_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__o32a_1
XFILLER_0_106_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24202_ clknet_leaf_117_clk _00735_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21414_ _03099_ _03097_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__and2b_1
X_22394_ _04066_ _04078_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24133_ clknet_leaf_0_clk _00666_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_21345_ _03076_ _03081_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__xor2_2
XFILLER_0_102_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_1123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24064_ clknet_leaf_83_clk _00597_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_21276_ _03013_ _03014_ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__nor2_1
XFILLER_0_241_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold650 top_inst.axis_out_inst.out_buff_data\[16\] VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 top_inst.axis_out_inst.out_buff_data\[23\] VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold672 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[31\] VGND
+ VGND VPWR VPWR net854 sky130_fd_sc_hd__dlygate4sd3_1
X_23015_ net33 net37 VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__nand2_2
Xhold683 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[23\] VGND
+ VGND VPWR VPWR net865 sky130_fd_sc_hd__dlygate4sd3_1
X_20227_ _02020_ _02021_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__or2_1
Xhold694 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[17\] VGND
+ VGND VPWR VPWR net876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20158_ _01968_ _01966_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__nand2_2
XFILLER_0_228_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12980_ _05748_ _05756_ _05769_ _05767_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__o211a_1
X_20089_ _01901_ _01902_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_239_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23917_ clknet_leaf_77_clk _00450_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ net665 _04969_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__or2_1
XTAP_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14650_ _07338_ _07339_ VGND VGND VPWR VPWR _07340_ sky130_fd_sc_hd__xor2_2
XTAP_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11862_ net367 _04930_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__or2_1
X_23848_ clknet_leaf_95_clk _00381_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13601_ _06306_ _06348_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _07256_ _07258_ VGND VGND VPWR VPWR _07272_ sky130_fd_sc_hd__or2_1
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23779_ clknet_leaf_65_clk _00312_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11793_ net829 _04885_ _04896_ _04889_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16320_ _08893_ _08849_ _08901_ VGND VGND VPWR VPWR _08902_ sky130_fd_sc_hd__o21a_1
XFILLER_0_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13532_ _06243_ _06256_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16251_ top_inst.grid_inst.data_path_wires\[8\]\[0\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _08834_ sky130_fd_sc_hd__or2b_1
XFILLER_0_137_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13463_ _05317_ _06217_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15202_ _07841_ _07797_ _07849_ VGND VGND VPWR VPWR _07850_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12414_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[22\] _05248_
+ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16182_ _08765_ _08766_ VGND VGND VPWR VPWR _08767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13394_ _05886_ _06166_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__and2_1
XFILLER_0_180_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15133_ top_inst.grid_inst.data_path_wires\[6\]\[0\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _07782_ sky130_fd_sc_hd__or2b_1
XFILLER_0_65_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12345_ net286 _05209_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1091 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19941_ _01395_ VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__buf_2
X_15064_ _07613_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[2\] _07712_
+ _07713_ VGND VGND VPWR VPWR _07715_ sky130_fd_sc_hd__nand4_2
XFILLER_0_239_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12276_ net906 _05164_ _05172_ _05168_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__o211a_1
X_14015_ _06364_ _06732_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19872_ _01671_ _01674_ _01694_ _10957_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__a31o_1
X_18823_ _11214_ _11215_ _11248_ VGND VGND VPWR VPWR _11249_ sky130_fd_sc_hd__a21o_1
XTAP_6160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18754_ _11171_ _11172_ VGND VGND VPWR VPWR _11183_ sky130_fd_sc_hd__nand2_1
X_15966_ _08568_ _08569_ _08575_ VGND VGND VPWR VPWR _08576_ sky130_fd_sc_hd__and3_1
XFILLER_0_234_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14917_ net229 _07597_ _07594_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__o21a_1
X_17705_ _10169_ _10214_ VGND VGND VPWR VPWR _10215_ sky130_fd_sc_hd__xnor2_1
XTAP_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18685_ _10577_ _10584_ _11131_ _10620_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15897_ _08478_ _08479_ _08508_ VGND VGND VPWR VPWR _08509_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_172_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_1004 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14848_ _07531_ _07528_ _07530_ VGND VGND VPWR VPWR _07533_ sky130_fd_sc_hd__or3_1
XFILLER_0_157_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17636_ _10099_ _10121_ _10147_ VGND VGND VPWR VPWR _10148_ sky130_fd_sc_hd__o21a_1
XFILLER_0_216_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17567_ _10069_ _10081_ VGND VGND VPWR VPWR _10082_ sky130_fd_sc_hd__xnor2_1
X_14779_ _07415_ _07465_ VGND VGND VPWR VPWR _07466_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19306_ top_inst.skew_buff_inst.row\[3\].output_reg\[6\] top_inst.axis_in_inst.inbuf_bus\[30\]
+ net188 VGND VGND VPWR VPWR _11704_ sky130_fd_sc_hd__mux2_4
X_16518_ _09055_ _09094_ VGND VGND VPWR VPWR _09095_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17498_ _10027_ _07611_ _10028_ _10024_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16449_ _09026_ _09027_ VGND VGND VPWR VPWR _09028_ sky130_fd_sc_hd__xnor2_1
X_19237_ _11645_ _11651_ VGND VGND VPWR VPWR _11652_ sky130_fd_sc_hd__xor2_1
XFILLER_0_147_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19168_ _11505_ _11543_ _11581_ _11584_ _11580_ VGND VGND VPWR VPWR _11585_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18119_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _10600_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19099_ _11516_ _11517_ VGND VGND VPWR VPWR _11518_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21130_ _02882_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21061_ _02824_ _02825_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__or2_1
X_20012_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[24\] _01764_ VGND
+ VGND VPWR VPWR _01829_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21963_ _03663_ _03664_ _03671_ _03676_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23702_ clknet_leaf_125_clk net601 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_20914_ _02684_ VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__clkbuf_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21894_ _03576_ _03596_ _03574_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23633_ clknet_leaf_103_clk _00166_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20845_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[20\] _02470_ VGND
+ VGND VPWR VPWR _02618_ sky130_fd_sc_hd__or2_1
XFILLER_0_232_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23564_ clknet_leaf_102_clk _00097_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20776_ _02549_ _02550_ _02466_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22515_ _04061_ _04195_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23495_ clknet_leaf_143_clk _00028_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[85\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22446_ _04061_ _04128_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22377_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[12\] _03894_ VGND
+ VGND VPWR VPWR _04062_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12130_ _05009_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__buf_2
XFILLER_0_66_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24116_ clknet_leaf_12_clk _00649_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_21328_ _03064_ _03065_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__nor2_1
XFILLER_0_237_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24047_ clknet_leaf_34_clk _00580_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_12061_ _05009_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__clkbuf_2
X_21259_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[5\] _02974_ _02975_
+ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_236_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold480 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[2\] VGND VGND
+ VPWR VPWR net662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold491 top_inst.axis_out_inst.out_buff_data\[33\] VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_216_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15820_ _08391_ _08396_ _08432_ _07439_ VGND VGND VPWR VPWR _08434_ sky130_fd_sc_hd__a31o_1
XFILLER_0_176_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_231_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15751_ _08360_ _08365_ VGND VGND VPWR VPWR _08366_ sky130_fd_sc_hd__xnor2_1
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12963_ _05757_ _05294_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__or2_1
XTAP_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_84_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _07387_ _07388_ _07371_ VGND VGND VPWR VPWR _07391_ sky130_fd_sc_hd__a21oi_1
XTAP_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11914_ net954 _04964_ _04965_ _04955_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18470_ _10853_ _10932_ VGND VGND VPWR VPWR _10933_ sky130_fd_sc_hd__xnor2_4
XTAP_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15682_ _08296_ _08297_ _08272_ _08273_ VGND VGND VPWR VPWR _08299_ sky130_fd_sc_hd__o211a_1
X_12894_ net998 _05403_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _09919_ _09957_ VGND VGND VPWR VPWR _09959_ sky130_fd_sc_hd__and2_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _07321_ _07320_ VGND VGND VPWR VPWR _07323_ sky130_fd_sc_hd__and2b_1
XFILLER_0_206_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11845_ net325 _04925_ _04926_ _04916_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__o211a_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _09871_ _09875_ _09874_ VGND VGND VPWR VPWR _09893_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14564_ _07253_ _07254_ _07255_ VGND VGND VPWR VPWR _07256_ sky130_fd_sc_hd__and3_1
XFILLER_0_173_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_947 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ top_inst.axis_out_inst.out_buff_data\[68\] _04877_ VGND VGND VPWR VPWR _04887_
+ sky130_fd_sc_hd__or2_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16303_ _08673_ _08693_ _08671_ _08690_ VGND VGND VPWR VPWR _08885_ sky130_fd_sc_hd__nand4_4
XFILLER_0_144_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13515_ top_inst.grid_inst.data_path_wires\[2\]\[1\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[2\]\[2\]
+ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__a22o_1
X_17283_ _09822_ _09827_ VGND VGND VPWR VPWR _09828_ sky130_fd_sc_hd__xnor2_1
X_14495_ _07161_ _07188_ VGND VGND VPWR VPWR _07189_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19022_ top_inst.grid_inst.data_path_wires\[13\]\[3\] top_inst.grid_inst.data_path_wires\[13\]\[4\]
+ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _11443_ sky130_fd_sc_hd__and4b_1
XFILLER_0_137_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16234_ _08815_ _08816_ _08817_ VGND VGND VPWR VPWR _08818_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13446_ _05260_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16165_ _08693_ _08690_ top_inst.grid_inst.data_path_wires\[8\]\[1\] top_inst.grid_inst.data_path_wires\[8\]\[0\]
+ VGND VGND VPWR VPWR _08751_ sky130_fd_sc_hd__nand4_1
XFILLER_0_106_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13377_ _06147_ _06148_ _06149_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_144_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15116_ _07719_ _07727_ VGND VGND VPWR VPWR _07766_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12328_ net319 _05196_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__or2_1
X_16096_ _08690_ _08684_ VGND VGND VPWR VPWR _08691_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19924_ _01743_ _01744_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__xor2_2
XFILLER_0_142_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15047_ _07696_ _07698_ VGND VGND VPWR VPWR _07699_ sky130_fd_sc_hd__xor2_2
X_12259_ net907 _05151_ _05162_ _05155_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19855_ _01657_ _01667_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__or2_1
XFILLER_0_235_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18806_ _11138_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[2\] VGND
+ VGND VPWR VPWR _11232_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19786_ _01604_ _01612_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_235_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16998_ _09549_ _09550_ _09465_ VGND VGND VPWR VPWR _09552_ sky130_fd_sc_hd__o21ai_4
X_18737_ _11149_ _11130_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _11168_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15949_ _08150_ _08353_ _08558_ VGND VGND VPWR VPWR _08559_ sky130_fd_sc_hd__o21a_1
XFILLER_0_183_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_75_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18668_ _11118_ _11124_ VGND VGND VPWR VPWR _11125_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_231_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17619_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[3\] _10129_ _10130_
+ VGND VGND VPWR VPWR _10131_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_231_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18599_ _11018_ _11021_ _11057_ VGND VGND VPWR VPWR _11059_ sky130_fd_sc_hd__and3_1
XFILLER_0_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20630_ _02403_ _02410_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_749 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20561_ _02269_ _02267_ _02307_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22300_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[5\] _03690_ VGND
+ VGND VPWR VPWR _03987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23280_ _04686_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__clkbuf_2
X_20492_ _01999_ _02015_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[9\]
+ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_950 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22231_ _03874_ _03849_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__or2b_1
XFILLER_0_162_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22162_ top_inst.grid_inst.data_path_wires\[18\]\[6\] top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[1\]
+ _03697_ _03695_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__a22o_1
XFILLER_0_219_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21113_ _01995_ _11142_ _02870_ _02707_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22093_ _03779_ _03784_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_1363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21044_ _02762_ _02805_ _02808_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__o21a_1
XFILLER_0_227_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22995_ net633 _04583_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_66_clk clknet_4_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21946_ top_inst.deskew_buff_inst.col_input\[94\] _03658_ _06140_ VGND VGND VPWR
+ VPWR _03661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21877_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[25\] _03421_ _03422_
+ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_167_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23616_ clknet_leaf_105_clk net539 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20828_ _02518_ _02601_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24596_ clknet_leaf_22_clk _01129_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23547_ clknet_leaf_103_clk net521 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20759_ _02486_ _02511_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__nor2_1
X_13300_ _06073_ _06075_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14280_ _06953_ _06955_ VGND VGND VPWR VPWR _06991_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23478_ clknet_leaf_134_clk net349 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13231_ top_inst.grid_inst.data_path_wires\[1\]\[3\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22429_ _04064_ _04065_ _04078_ _04077_ _04075_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__o32a_1
XFILLER_0_126_1015 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13162_ _05894_ _05897_ _05898_ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_1183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12113_ net262 _05071_ _05079_ _05075_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13093_ _05849_ _05850_ _05873_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__a21oi_1
X_17970_ _10430_ _10432_ VGND VGND VPWR VPWR _10474_ sky130_fd_sc_hd__or2b_1
XFILLER_0_27_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16921_ _09473_ _09474_ _09475_ VGND VGND VPWR VPWR _09477_ sky130_fd_sc_hd__a21o_1
X_12044_ net264 _05036_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__or2_1
XFILLER_0_178_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19640_ _01467_ _01469_ _05399_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__a21oi_1
X_16852_ _09402_ _09404_ _09401_ VGND VGND VPWR VPWR _09409_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_244_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_217_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15803_ _08362_ _08364_ _08416_ VGND VGND VPWR VPWR _08417_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_232_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16783_ _09308_ _09340_ _09341_ VGND VGND VPWR VPWR _09342_ sky130_fd_sc_hd__nand3_2
X_19571_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[3\]
+ _11700_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__and3_1
XFILLER_0_189_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13995_ _06711_ _06712_ VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_57_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_233_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15734_ _08342_ _08343_ _08348_ VGND VGND VPWR VPWR _08349_ sky130_fd_sc_hd__a21o_1
X_18522_ _10933_ _10983_ VGND VGND VPWR VPWR _10984_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12946_ _05744_ _05735_ _05745_ _05743_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__o211a_1
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15665_ _08276_ _08281_ VGND VGND VPWR VPWR _08282_ sky130_fd_sc_hd__xnor2_1
X_18453_ _10881_ _10916_ VGND VGND VPWR VPWR _10917_ sky130_fd_sc_hd__nand2_1
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12877_ _05608_ _05649_ _05647_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__a21o_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17404_ _09911_ _09921_ _09938_ _09899_ VGND VGND VPWR VPWR _09943_ sky130_fd_sc_hd__a22o_1
X_14616_ _07261_ _07263_ VGND VGND VPWR VPWR _07307_ sky130_fd_sc_hd__nand2_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11828_ _04876_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__buf_2
X_18384_ top_inst.grid_inst.data_path_wires\[12\]\[5\] _10608_ _10604_ _10591_ VGND
+ VGND VPWR VPWR _10849_ sky130_fd_sc_hd__a22o_1
X_15596_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[3\] _05326_ VGND
+ VGND VPWR VPWR _08216_ sky130_fd_sc_hd__and2_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17335_ _09854_ _09876_ VGND VGND VPWR VPWR _09877_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _07237_ _07238_ VGND VGND VPWR VPWR _07239_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11759_ top_inst.axis_out_inst.out_buff_data\[124\] _04877_ VGND VGND VPWR VPWR _04878_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_12_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17266_ _09625_ _09793_ VGND VGND VPWR VPWR _09811_ sky130_fd_sc_hd__nor2_1
X_14478_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[3\]
+ _07064_ _07068_ VGND VGND VPWR VPWR _07172_ sky130_fd_sc_hd__nand4_4
XFILLER_0_181_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16217_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[3\]
+ top_inst.grid_inst.data_path_wires\[8\]\[3\] _08667_ VGND VGND VPWR VPWR _08801_
+ sky130_fd_sc_hd__nand4_2
X_19005_ _11375_ _11377_ _11422_ VGND VGND VPWR VPWR _11426_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13429_ _05748_ _06192_ _06194_ _06183_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17197_ _09744_ _09745_ VGND VGND VPWR VPWR _09746_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16148_ _08727_ _08734_ VGND VGND VPWR VPWR _08735_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16079_ _08150_ _08663_ _08678_ _08666_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19907_ _01720_ _01728_ VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_227_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_243_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19838_ _01658_ _01661_ _01662_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__nand3_1
XFILLER_0_224_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_235_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 input_tdata[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_4
X_19769_ _01588_ _01589_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__or2b_1
Xclkbuf_leaf_48_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_155_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21800_ _03503_ _03521_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22780_ _04192_ _04431_ _04448_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__nand3_1
XFILLER_0_91_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21731_ _03446_ _03455_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24450_ clknet_leaf_64_clk _00983_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21662_ _03389_ _03390_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23401_ net64 _04658_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20613_ _02356_ _02359_ net174 _02393_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__o31a_1
X_24381_ clknet_leaf_38_clk _00914_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21593_ _03287_ _03288_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23332_ net157 _04779_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20544_ _02325_ _02326_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__xor2_1
XFILLER_0_132_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23263_ net124 _04740_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20475_ _02222_ _02259_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22214_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[5\] _03686_ VGND
+ VGND VPWR VPWR _03903_ sky130_fd_sc_hd__nand2_1
X_23194_ net91 _04701_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22145_ _03809_ _03810_ _03834_ _03835_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_24_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22076_ _03765_ _03768_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__xor2_2
XTAP_6759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21027_ _02643_ _02792_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__xor2_2
XFILLER_0_227_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_214_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_39_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_199_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12800_ _05606_ _05607_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__nor2_2
XFILLER_0_214_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13780_ _06491_ _06490_ VGND VGND VPWR VPWR _06523_ sky130_fd_sc_hd__or2b_1
X_22978_ net633 _04575_ _04579_ _04577_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12731_ _05534_ _05539_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21929_ _03622_ _03640_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15450_ _08058_ _08091_ VGND VGND VPWR VPWR _08092_ sky130_fd_sc_hd__nor2_1
X_12662_ _05443_ _05429_ _05472_ _05473_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14401_ _07096_ _07097_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[1\]
+ VGND VGND VPWR VPWR _07099_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15381_ _08022_ _08024_ VGND VGND VPWR VPWR _08025_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24579_ clknet_leaf_140_clk _01112_ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dfxtp_4
X_12593_ _05405_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__buf_8
XFILLER_0_93_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17120_ _09553_ _09641_ _09640_ VGND VGND VPWR VPWR _09671_ sky130_fd_sc_hd__o21ba_1
X_14332_ _07039_ _07040_ VGND VGND VPWR VPWR _07041_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17051_ _09553_ _09602_ _09603_ VGND VGND VPWR VPWR _09604_ sky130_fd_sc_hd__or3_1
XFILLER_0_145_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_1304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14263_ _06961_ _06962_ _06973_ VGND VGND VPWR VPWR _06974_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16002_ _08593_ _08576_ _08609_ VGND VGND VPWR VPWR _08611_ sky130_fd_sc_hd__or3_1
X_13214_ _05986_ _05991_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__xnor2_1
X_14194_ _06825_ _06906_ VGND VGND VPWR VPWR _06907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_237_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13145_ _05924_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13076_ top_inst.grid_inst.data_path_wires\[1\]\[2\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[1\]\[3\]
+ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__a22o_1
X_17953_ _10452_ _10456_ VGND VGND VPWR VPWR _10457_ sky130_fd_sc_hd__xnor2_2
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16904_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[8\] _09459_ _09417_
+ VGND VGND VPWR VPWR _09460_ sky130_fd_sc_hd__a21o_1
X_12027_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[16\] _05023_
+ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__or2_1
X_17884_ _10387_ _10389_ VGND VGND VPWR VPWR _10390_ sky130_fd_sc_hd__xor2_1
XFILLER_0_228_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19623_ _01451_ _01452_ _01444_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__a21o_1
XFILLER_0_217_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16835_ _09329_ _09331_ _09391_ _09392_ VGND VGND VPWR VPWR _09393_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19554_ net846 _01386_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__or2_1
XFILLER_0_233_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16766_ _09193_ _09209_ _09214_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _09325_ sky130_fd_sc_hd__a22o_1
X_13978_ _06676_ _06696_ VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18505_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[11\] _10923_ _10840_
+ VGND VGND VPWR VPWR _10967_ sky130_fd_sc_hd__a21o_1
XFILLER_0_232_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12929_ _05715_ _05719_ _05729_ _05732_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__a31o_1
XFILLER_0_186_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15717_ _08323_ _08332_ VGND VGND VPWR VPWR _08333_ sky130_fd_sc_hd__xor2_1
X_16697_ _09258_ VGND VGND VPWR VPWR _09259_ sky130_fd_sc_hd__inv_2
X_19485_ _01275_ _01317_ _01318_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__nand3_1
XFILLER_0_220_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18436_ _10896_ _10899_ VGND VGND VPWR VPWR _10900_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15648_ _08237_ _08263_ _08265_ VGND VGND VPWR VPWR _08266_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18367_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[8\] _09496_ _10830_
+ _10832_ VGND VGND VPWR VPWR _10833_ sky130_fd_sc_hd__a22o_1
X_15579_ _08135_ _08161_ _08159_ _08137_ VGND VGND VPWR VPWR _08199_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17318_ _09844_ _09860_ VGND VGND VPWR VPWR _09861_ sky130_fd_sc_hd__or2_1
XFILLER_0_173_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18298_ _10589_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[2\] _10762_
+ _10763_ VGND VGND VPWR VPWR _10765_ sky130_fd_sc_hd__nand4_1
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17249_ _09792_ _09794_ VGND VGND VPWR VPWR _09795_ sky130_fd_sc_hd__xor2_2
XFILLER_0_189_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20260_ _02030_ _02044_ _02045_ VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__or3b_1
XFILLER_0_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20191_ _01995_ _10033_ _01996_ _01840_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__o211a_1
XFILLER_0_228_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23950_ clknet_leaf_90_clk _00483_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22901_ _10583_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__clkbuf_4
XTAP_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23881_ clknet_leaf_50_clk _00414_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22832_ _10583_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22763_ _04432_ _04431_ _04412_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24502_ clknet_leaf_123_clk _01035_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_220_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21714_ _03399_ _03439_ _03440_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_91_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22694_ _04331_ _04366_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__and2_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24433_ clknet_leaf_57_clk net607 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_21645_ _03210_ _03328_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__and2b_1
XFILLER_0_240_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24364_ clknet_leaf_31_clk _00897_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[123\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_50 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21576_ _03269_ _03307_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__xnor2_1
XANTENNA_61 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_72 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23315_ net149 _04766_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__or2_1
XANTENNA_83 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20527_ net883 _01735_ _02310_ _02035_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_94 net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24295_ clknet_leaf_137_clk _00828_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23246_ net116 _04727_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20458_ top_inst.grid_inst.data_path_wires\[16\]\[6\] top_inst.grid_inst.data_path_wires\[16\]\[5\]
+ _02013_ _02011_ VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__nand4_1
XFILLER_0_132_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23177_ net83 _04687_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__or2_1
XTAP_6501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20389_ _02129_ _02127_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_242_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22128_ _03813_ _03818_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__xor2_1
XTAP_6534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14950_ _07617_ VGND VGND VPWR VPWR _07618_ sky130_fd_sc_hd__buf_2
X_22059_ _03737_ _03751_ _03752_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__nand3_1
XTAP_6589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13901_ _06196_ _06192_ _06633_ _06446_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__o211a_1
X_14881_ _07532_ _07564_ VGND VGND VPWR VPWR _07565_ sky130_fd_sc_hd__xor2_1
XTAP_5888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16620_ net1119 VGND VGND VPWR VPWR _09192_ sky130_fd_sc_hd__clkbuf_4
X_13832_ _06572_ _06573_ VGND VGND VPWR VPWR _06574_ sky130_fd_sc_hd__nor2_1
XFILLER_0_216_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_1125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16551_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[14\] _08975_ VGND
+ VGND VPWR VPWR _09127_ sky130_fd_sc_hd__xnor2_1
X_13763_ _06385_ _06506_ VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_1135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12714_ _05483_ _05524_ _05440_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__a21oi_1
X_15502_ top_inst.grid_inst.data_path_wires\[7\]\[2\] VGND VGND VPWR VPWR _08139_
+ sky130_fd_sc_hd__clkbuf_4
X_16482_ _09054_ _09059_ VGND VGND VPWR VPWR _09060_ sky130_fd_sc_hd__xnor2_2
X_19270_ net1032 _11662_ _11675_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__o21a_1
XFILLER_0_195_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13694_ _06393_ _06395_ VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15433_ _08068_ _08038_ _08073_ VGND VGND VPWR VPWR _08075_ sky130_fd_sc_hd__nand3_1
XFILLER_0_127_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18221_ _10684_ _10689_ VGND VGND VPWR VPWR _10690_ sky130_fd_sc_hd__xnor2_2
X_12645_ _05455_ _05456_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__or2_1
XFILLER_0_182_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15364_ _08005_ _08006_ VGND VGND VPWR VPWR _08008_ sky130_fd_sc_hd__and2_1
X_18152_ _10623_ _10624_ _10617_ VGND VGND VPWR VPWR _10625_ sky130_fd_sc_hd__a21o_1
X_12576_ _05383_ _05389_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17103_ _09587_ _09613_ VGND VGND VPWR VPWR _09655_ sky130_fd_sc_hd__nand2_1
X_14315_ _07024_ VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18083_ net639 _10563_ _10576_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15295_ _07939_ _07940_ VGND VGND VPWR VPWR _07941_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17034_ _09544_ _09547_ _09586_ VGND VGND VPWR VPWR _09587_ sky130_fd_sc_hd__a21o_1
X_14246_ _06956_ _06957_ VGND VGND VPWR VPWR _06958_ sky130_fd_sc_hd__xnor2_1
Xhold309 _00230_ VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14177_ top_inst.grid_inst.data_path_wires\[3\]\[3\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _06890_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _05906_ _05907_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__or2_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18985_ _11161_ _11138_ _11352_ _11350_ VGND VGND VPWR VPWR _11407_ sky130_fd_sc_hd__a31oi_2
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _05802_ _05815_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__nand2_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17936_ _10439_ _10440_ VGND VGND VPWR VPWR _10441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17867_ _10371_ _10372_ VGND VGND VPWR VPWR _10373_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19606_ _11688_ _11709_ _01404_ _01403_ _11705_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__a32o_1
X_16818_ _09211_ _09197_ VGND VGND VPWR VPWR _09376_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17798_ _10297_ _10305_ VGND VGND VPWR VPWR _10306_ sky130_fd_sc_hd__xor2_1
XFILLER_0_117_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19537_ _01366_ _01367_ _01368_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__a21o_1
X_16749_ _09211_ _09187_ _09306_ _09307_ VGND VGND VPWR VPWR _09309_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_177_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19468_ _11683_ _11704_ _11708_ _11678_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18419_ _10870_ _10839_ VGND VGND VPWR VPWR _10883_ sky130_fd_sc_hd__or2b_1
XFILLER_0_185_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19399_ _01232_ _01233_ _01213_ _01215_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_5_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21430_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[10\] _03080_ VGND
+ VGND VPWR VPWR _03165_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_228_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21361_ _03009_ _03054_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23100_ net605 _10541_ _04648_ _04643_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20312_ _02086_ _02087_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__nand2_1
X_24080_ clknet_leaf_113_clk _00613_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold810 top_inst.axis_in_inst.inbuf_bus\[9\] VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21292_ top_inst.deskew_buff_inst.col_input\[70\] _03030_ _06140_ VGND VGND VPWR
+ VPWR _03031_ sky130_fd_sc_hd__mux2_1
Xhold821 top_inst.axis_in_inst.inbuf_bus\[30\] VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 top_inst.deskew_buff_inst.col_input\[96\] VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__dlymetal6s2s_1
X_23031_ net28 _04601_ _04610_ _04606_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold843 top_inst.axis_out_inst.out_buff_data\[58\] VGND VGND VPWR VPWR net1025 sky130_fd_sc_hd__dlygate4sd3_1
X_20243_ _10447_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold854 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[2\] VGND VGND
+ VPWR VPWR net1036 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold865 top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[23\] VGND VGND
+ VPWR VPWR net1047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR net1058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 _00532_ VGND VGND VPWR VPWR net1069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold898 top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[16\] VGND VGND
+ VPWR VPWR net1080 sky130_fd_sc_hd__dlygate4sd3_1
X_20174_ _05633_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__buf_8
XTAP_5107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1062 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23933_ clknet_leaf_85_clk _00466_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_157_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23864_ clknet_leaf_68_clk _00397_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22815_ _04444_ _04480_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_233_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23795_ clknet_leaf_69_clk _00328_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_39_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22746_ _04415_ _04416_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__nand2_1
XFILLER_0_177_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22677_ _04349_ _04350_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24416_ clknet_leaf_56_clk _00949_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12430_ _04868_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21628_ _03356_ _03357_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_1287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24347_ clknet_leaf_26_clk _00880_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[106\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12361_ _05127_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21559_ _03254_ _03255_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__or2b_1
X_14100_ _06648_ top_inst.grid_inst.data_path_wires\[3\]\[4\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[3\]
+ top_inst.grid_inst.data_path_wires\[3\]\[5\] VGND VGND VPWR VPWR _06815_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15080_ _07693_ _07694_ _07730_ VGND VGND VPWR VPWR _07731_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12292_ _05127_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__buf_2
X_24278_ clknet_leaf_12_clk _00811_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[17\]\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_105_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14031_ _06742_ _06747_ VGND VGND VPWR VPWR _06748_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_142_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23229_ net108 _04714_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18770_ _11195_ _11196_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[3\]
+ VGND VGND VPWR VPWR _11198_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15982_ _08588_ _08590_ _08591_ VGND VGND VPWR VPWR _08592_ sky130_fd_sc_hd__o21ai_1
XTAP_6386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17721_ _10197_ _10201_ VGND VGND VPWR VPWR _10230_ sky130_fd_sc_hd__nor2_1
X_14933_ _07592_ _07605_ _04870_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__o21a_1
XTAP_5674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ _10161_ _10162_ VGND VGND VPWR VPWR _10163_ sky130_fd_sc_hd__nand2_1
X_14864_ _07514_ _07547_ VGND VGND VPWR VPWR _07549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16603_ _09055_ _09153_ _09176_ VGND VGND VPWR VPWR _09177_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13815_ top_inst.grid_inst.data_path_wires\[2\]\[7\] _06214_ VGND VGND VPWR VPWR
+ _06557_ sky130_fd_sc_hd__nand2_1
X_14795_ _07480_ _07481_ _06682_ VGND VGND VPWR VPWR _07482_ sky130_fd_sc_hd__a21o_1
XFILLER_0_187_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17583_ _10095_ _10096_ VGND VGND VPWR VPWR _10097_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19322_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[1\] _11715_ _11716_
+ VGND VGND VPWR VPWR _11717_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16534_ _09069_ _09110_ VGND VGND VPWR VPWR _09111_ sky130_fd_sc_hd__xor2_1
X_13746_ _06488_ _06489_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19253_ _11646_ _11650_ VGND VGND VPWR VPWR _11667_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16465_ _08697_ _08676_ _09041_ VGND VGND VPWR VPWR _09043_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13677_ _06417_ _06422_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18204_ _10671_ _10673_ VGND VGND VPWR VPWR _10674_ sky130_fd_sc_hd__xor2_2
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12628_ _05404_ _05439_ _05440_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15416_ _08055_ _08057_ VGND VGND VPWR VPWR _08059_ sky130_fd_sc_hd__or2_1
X_16396_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[9\] _08975_ _08896_
+ VGND VGND VPWR VPWR _08976_ sky130_fd_sc_hd__a21o_1
X_19184_ _11597_ _11600_ VGND VGND VPWR VPWR _11601_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15347_ _07619_ _07824_ VGND VGND VPWR VPWR _07991_ sky130_fd_sc_hd__nor2_1
X_18135_ _10589_ _10607_ _10611_ _10594_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12559_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[4\] _05354_ _05372_
+ _05373_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15278_ _07845_ VGND VGND VPWR VPWR _07924_ sky130_fd_sc_hd__clkbuf_4
X_18066_ _10413_ _10549_ _10548_ VGND VGND VPWR VPWR _10566_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold106 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[26\] VGND
+ VGND VPWR VPWR net288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold117 _00284_ VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold128 top_inst.axis_out_inst.out_buff_data\[8\] VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17017_ _09542_ _09569_ _09570_ VGND VGND VPWR VPWR _09571_ sky130_fd_sc_hd__and3_1
X_14229_ _06937_ _06940_ VGND VGND VPWR VPWR _06941_ sky130_fd_sc_hd__nor2_1
Xhold139 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[23\] VGND
+ VGND VPWR VPWR net321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_226_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18968_ _11345_ _11347_ _11389_ VGND VGND VPWR VPWR _11390_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_193_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17919_ _10421_ _10422_ _10419_ VGND VGND VPWR VPWR _10424_ sky130_fd_sc_hd__o21a_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18899_ _11299_ _11322_ VGND VGND VPWR VPWR _11323_ sky130_fd_sc_hd__xor2_1
XFILLER_0_217_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20930_ _02698_ _02699_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__and2_1
XFILLER_0_179_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20861_ _02586_ _02593_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__nor2_1
X_22600_ _04248_ _04277_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23580_ clknet_leaf_106_clk _00113_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_20792_ net280 _02491_ _02566_ _02567_ _01863_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__o221a_1
XFILLER_0_152_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22531_ _04210_ _04188_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__or2b_1
XFILLER_0_14_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22462_ _04132_ _04144_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24201_ clknet_leaf_116_clk _00734_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21413_ _03130_ _03148_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_162_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22393_ _04075_ _04077_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24132_ clknet_leaf_4_clk _00665_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_21344_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[8\] _03080_ VGND
+ VGND VPWR VPWR _03081_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24063_ clknet_leaf_83_clk _00596_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold640 top_inst.axis_out_inst.out_buff_data\[41\] VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21275_ _02871_ _02887_ _03011_ _03012_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__o2bb2a_1
Xhold651 top_inst.axis_out_inst.out_buff_data\[108\] VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold662 top_inst.axis_out_inst.out_buff_data\[35\] VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__dlygate4sd3_1
X_23014_ net258 _04588_ _04599_ _04590_ VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold673 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[12\] VGND
+ VGND VPWR VPWR net855 sky130_fd_sc_hd__dlygate4sd3_1
X_20226_ _05772_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_229_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold684 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[10\] VGND
+ VGND VPWR VPWR net866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_228_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold695 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[0\] VGND
+ VGND VPWR VPWR net877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20157_ _01912_ _01929_ _01947_ _01967_ _01946_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__a32o_2
XFILLER_0_243_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_239_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20088_ _01870_ _01877_ _01897_ _01850_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__a22oi_2
XTAP_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ net970 _04964_ _04974_ _04968_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__o211a_1
X_23916_ clknet_leaf_35_clk _00449_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11861_ net808 _04925_ _04935_ _04929_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__o211a_1
X_23847_ clknet_leaf_95_clk _00380_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _06341_ _06347_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14580_ _07271_ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23778_ clknet_leaf_64_clk _00311_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11792_ net727 _04890_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13531_ _06279_ _06280_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__xor2_1
X_22729_ _04398_ _04400_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16250_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[8\]\[1\]
+ VGND VGND VPWR VPWR _08833_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13462_ _06181_ _06200_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15201_ _07847_ _07848_ VGND VGND VPWR VPWR _07849_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12413_ net298 _05243_ _05250_ _05247_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16181_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[3\]
+ _08667_ top_inst.grid_inst.data_path_wires\[8\]\[1\] VGND VGND VPWR VPWR _08766_
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13393_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[14\] _05354_ _06164_
+ _06165_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15132_ top_inst.grid_inst.data_path_wires\[6\]\[1\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _07781_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12344_ net726 _05204_ _05211_ _05208_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_239_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19940_ _01738_ _01742_ _01740_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__a21o_1
X_15063_ _07613_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[2\] _07712_
+ _07713_ VGND VGND VPWR VPWR _07714_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12275_ net747 _05169_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__or2_1
XFILLER_0_181_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14014_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[5\] _06242_ _06730_
+ _06731_ VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19871_ _01671_ _01674_ _01694_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__a21oi_1
X_18822_ _11193_ _11213_ VGND VGND VPWR VPWR _11248_ sky130_fd_sc_hd__nor2_1
XTAP_6150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18753_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[2\] _11181_ VGND
+ VGND VPWR VPWR _11182_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_218_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15965_ _08570_ _08574_ VGND VGND VPWR VPWR _08575_ sky130_fd_sc_hd__xor2_1
XTAP_5471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17704_ _10210_ _10213_ VGND VGND VPWR VPWR _10214_ sky130_fd_sc_hd__xnor2_1
X_14916_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[18\] _07595_ VGND
+ VGND VPWR VPWR _07597_ sky130_fd_sc_hd__and2_1
XTAP_5493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18684_ _11130_ _08674_ VGND VGND VPWR VPWR _11131_ sky130_fd_sc_hd__or2_1
XFILLER_0_236_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15896_ _08505_ _08507_ VGND VGND VPWR VPWR _08508_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_215_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1016 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17635_ _10118_ _10120_ VGND VGND VPWR VPWR _10147_ sky130_fd_sc_hd__or2b_1
X_14847_ _07528_ _07530_ _07531_ VGND VGND VPWR VPWR _07532_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17566_ _10079_ _10080_ VGND VGND VPWR VPWR _10081_ sky130_fd_sc_hd__and2_1
X_14778_ _07458_ _07464_ VGND VGND VPWR VPWR _07465_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19305_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _11703_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16517_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[13\] _08975_ VGND
+ VGND VPWR VPWR _09094_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13729_ _06430_ _06473_ VGND VGND VPWR VPWR _06474_ sky130_fd_sc_hd__xnor2_1
X_17497_ _05736_ _09197_ VGND VGND VPWR VPWR _10028_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19236_ _11646_ _11650_ VGND VGND VPWR VPWR _11651_ sky130_fd_sc_hd__xor2_1
XFILLER_0_171_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16448_ _08974_ _08980_ _08972_ VGND VGND VPWR VPWR _09027_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19167_ _11549_ _11548_ VGND VGND VPWR VPWR _11584_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16379_ _08927_ _08933_ _08958_ VGND VGND VPWR VPWR _08959_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18118_ top_inst.grid_inst.data_path_wires\[12\]\[1\] VGND VGND VPWR VPWR _10599_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19098_ _11513_ _11515_ VGND VGND VPWR VPWR _11517_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18049_ _10413_ _10549_ VGND VGND VPWR VPWR _10550_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21060_ _02810_ _02823_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20011_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[23\] _01761_ _01762_
+ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21962_ _03674_ _03675_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_193_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23701_ clknet_leaf_125_clk _00234_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20913_ _02135_ _02683_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__and2_1
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21893_ _03603_ _03604_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__or2b_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_230_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23632_ clknet_leaf_103_clk _00165_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20844_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[20\] _02468_ VGND
+ VGND VPWR VPWR _02617_ sky130_fd_sc_hd__nand2_1
XFILLER_0_230_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23563_ clknet_leaf_100_clk net792 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20775_ _02465_ _02549_ _02550_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22514_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[16\] _03894_ VGND
+ VGND VPWR VPWR _04195_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23494_ clknet_leaf_143_clk _00027_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[84\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22445_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[14\] _03894_ VGND
+ VGND VPWR VPWR _04128_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22376_ _04060_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_241_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24115_ clknet_leaf_118_clk _00648_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21327_ _03027_ _03029_ _03026_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_60_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_4__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_4_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_241_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24046_ clknet_4_7__leaf_clk _00579_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_12060_ net327 _05045_ _05048_ _05049_ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold470 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[25\] VGND
+ VGND VPWR VPWR net652 sky130_fd_sc_hd__dlygate4sd3_1
X_21258_ _02971_ _02979_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__and2_1
XFILLER_0_241_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold481 _00952_ VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold492 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[5\] VGND VGND
+ VPWR VPWR net674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20209_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _02009_ sky130_fd_sc_hd__clkbuf_4
X_21189_ _02928_ _02929_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[3\]
+ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_1152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12962_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _05757_ sky130_fd_sc_hd__clkbuf_4
XTAP_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _08363_ _08364_ VGND VGND VPWR VPWR _08365_ sky130_fd_sc_hd__nand2_1
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ _07389_ VGND VGND VPWR VPWR _07390_ sky130_fd_sc_hd__inv_2
XTAP_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ net428 _04956_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12893_ _05698_ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__clkbuf_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15681_ _08272_ _08273_ _08296_ _08297_ VGND VGND VPWR VPWR _08298_ sky130_fd_sc_hd__a211oi_2
XTAP_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17420_ _09919_ _09957_ VGND VGND VPWR VPWR _09958_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _07320_ _07321_ VGND VGND VPWR VPWR _07322_ sky130_fd_sc_hd__and2b_1
X_11844_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[1\] _04917_
+ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__or2_1
XTAP_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14563_ _07209_ _07211_ VGND VGND VPWR VPWR _07255_ sky130_fd_sc_hd__nand2_1
X_17351_ _09721_ _09824_ _09888_ _09891_ VGND VGND VPWR VPWR _09892_ sky130_fd_sc_hd__o31ai_4
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11775_ net594 _04885_ _04886_ _04875_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_200_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16302_ _08693_ _08671_ _08690_ _08673_ VGND VGND VPWR VPWR _08884_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_1370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ _06181_ _06212_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__nand2_1
X_17282_ _09721_ _09824_ _09826_ VGND VGND VPWR VPWR _09827_ sky130_fd_sc_hd__o21bai_2
X_14494_ _07185_ _07187_ VGND VGND VPWR VPWR _07188_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19021_ _11161_ _11143_ VGND VGND VPWR VPWR _11442_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16233_ _08770_ _08778_ VGND VGND VPWR VPWR _08817_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13445_ _06205_ _05773_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16164_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[2\] _08667_ VGND
+ VGND VPWR VPWR _08750_ sky130_fd_sc_hd__nand2_1
X_13376_ _05753_ _06082_ _06085_ _06115_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15115_ _07754_ _07763_ VGND VGND VPWR VPWR _07765_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12327_ net890 _05191_ _05201_ _05195_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__o211a_1
X_16095_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _08690_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19923_ _01611_ _01726_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__nor2_1
X_15046_ _07635_ _07670_ _07697_ VGND VGND VPWR VPWR _07698_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_220_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12258_ net863 _05156_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19854_ _01669_ _01654_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__or2b_1
X_12189_ top_inst.axis_out_inst.out_buff_data\[22\] _05115_ VGND VGND VPWR VPWR _05122_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_208_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18805_ _11161_ _11130_ VGND VGND VPWR VPWR _11231_ sky130_fd_sc_hd__nand2_1
X_19785_ _01606_ _01609_ _01610_ _01611_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__a211o_1
X_16997_ _09465_ _09549_ _09550_ VGND VGND VPWR VPWR _09551_ sky130_fd_sc_hd__or3_4
XFILLER_0_223_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18736_ _11149_ _11130_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _11167_ sky130_fd_sc_hd__and3_1
XTAP_5290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15948_ _08152_ _08169_ VGND VGND VPWR VPWR _08558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18667_ _11120_ _11123_ VGND VGND VPWR VPWR _11124_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15879_ _08489_ _08490_ VGND VGND VPWR VPWR _08491_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_203_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_231_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17618_ top_inst.grid_inst.data_path_wires\[11\]\[1\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[11\]\[2\]
+ VGND VGND VPWR VPWR _10130_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18598_ _11018_ _11021_ _11057_ VGND VGND VPWR VPWR _11058_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_231_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17549_ _10025_ _10022_ _10044_ _10042_ VGND VGND VPWR VPWR _10065_ sky130_fd_sc_hd__nand4_2
XFILLER_0_4_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20560_ _02311_ _02342_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__xor2_2
XFILLER_0_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19219_ _11633_ _11634_ VGND VGND VPWR VPWR _11635_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_1387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20491_ _01993_ _02227_ _02238_ _02239_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_144_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22230_ _03888_ _03918_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__xor2_2
XFILLER_0_229_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22161_ _03826_ _03827_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21112_ _02868_ _02869_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__or2_1
X_22092_ _03780_ _03783_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__xor2_2
XFILLER_0_26_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21043_ _02774_ _02778_ _02800_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_199_1375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_236_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22994_ _05736_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_4_12__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_4_12__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_242_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21945_ _03070_ _03658_ _03659_ _03660_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21876_ _03549_ _03593_ _03594_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_171_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23615_ clknet_leaf_105_clk net273 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20827_ _02574_ _02600_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__xnor2_1
X_24595_ clknet_leaf_23_clk _01128_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_166_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23546_ clknet_leaf_129_clk _00079_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20758_ _02508_ _02534_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23477_ clknet_leaf_136_clk _00010_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20689_ _02467_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__clkbuf_4
X_13230_ _05976_ _05981_ _06006_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22428_ _04099_ _04111_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__xor2_1
XFILLER_0_122_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13161_ _05934_ _05939_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__xnor2_1
X_22359_ _04042_ _04044_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__xor2_2
XFILLER_0_33_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12112_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[20\] _05076_
+ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_1363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13092_ _05852_ _05872_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16920_ _09473_ _09474_ _09475_ VGND VGND VPWR VPWR _09476_ sky130_fd_sc_hd__nand3_1
X_24029_ clknet_leaf_48_clk _00562_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12043_ net672 _05031_ _05039_ _05035_ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16851_ _09408_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_232_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15802_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[9\] _08374_ VGND
+ VGND VPWR VPWR _08416_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_219_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_217_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19570_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[2\] _11708_ VGND
+ VGND VPWR VPWR _01402_ sky130_fd_sc_hd__nand2_4
X_16782_ _09335_ _09336_ _09339_ VGND VGND VPWR VPWR _09341_ sky130_fd_sc_hd__a21o_1
XFILLER_0_176_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_232_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13994_ _06626_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[2\] _06709_
+ _06710_ VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__and4_1
X_18521_ _10981_ _10982_ VGND VGND VPWR VPWR _10983_ sky130_fd_sc_hd__xnor2_1
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ _08300_ _08341_ VGND VGND VPWR VPWR _08348_ sky130_fd_sc_hd__nor2_1
X_12945_ _05739_ _05528_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__nand2_1
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18452_ _10914_ _10915_ VGND VGND VPWR VPWR _10916_ sky130_fd_sc_hd__and2_1
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _08279_ _08280_ VGND VGND VPWR VPWR _08281_ sky130_fd_sc_hd__nand2_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12876_ _05680_ _05681_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17403_ _09940_ _09941_ VGND VGND VPWR VPWR _09942_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14615_ _07272_ _07305_ VGND VGND VPWR VPWR _07306_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ net652 _04912_ _04915_ _04916_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__o211a_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _10801_ _10809_ VGND VGND VPWR VPWR _10848_ sky130_fd_sc_hd__or2b_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15595_ _08212_ _08213_ _08195_ VGND VGND VPWR VPWR _08215_ sky130_fd_sc_hd__o21ai_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _09874_ _09875_ VGND VGND VPWR VPWR _09876_ sky130_fd_sc_hd__and2b_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14546_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[3\]
+ _07072_ _07077_ VGND VGND VPWR VPWR _07238_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11758_ _04876_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__buf_4
XFILLER_0_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17265_ _09774_ _09809_ VGND VGND VPWR VPWR _09810_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14477_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[4\] _07064_ _07068_
+ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _07171_ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19004_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[9\] _10364_ _11424_
+ _11425_ _11228_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__o221a_1
XFILLER_0_10_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16216_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[8\]\[3\]
+ _08667_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _08800_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13428_ _06193_ _05262_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17196_ _09721_ _09743_ VGND VGND VPWR VPWR _09745_ sky130_fd_sc_hd__nand2_1
XFILLER_0_178_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16147_ _08732_ _08733_ VGND VGND VPWR VPWR _08734_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_141_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13359_ _06113_ _06132_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16078_ _08677_ _08674_ VGND VGND VPWR VPWR _08678_ sky130_fd_sc_hd__or2_1
XFILLER_0_220_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19906_ _01726_ _01727_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__xor2_2
X_15029_ _07681_ VGND VGND VPWR VPWR _07682_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19837_ _01659_ _01660_ _01528_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_242_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19768_ _01518_ _01556_ _01591_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__nor3_1
Xinput2 input_tdata[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_4
XFILLER_0_155_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18719_ _11135_ _10607_ _11155_ _11137_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19699_ _01527_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__buf_4
XFILLER_0_151_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21730_ _03446_ _03455_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_210_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21661_ _03387_ _03388_ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_231_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23400_ net451 _04655_ _04820_ _04819_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20612_ _02355_ _02362_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__or2b_1
X_24380_ clknet_leaf_39_clk _00913_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1054 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21592_ _03287_ _03288_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23331_ net599 _04778_ _04781_ _04782_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20543_ _01999_ _02018_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23262_ net1059 _04739_ _04742_ _04743_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20474_ _02257_ _02258_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22213_ _03900_ _03901_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23193_ net972 _04700_ _04703_ _04704_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22144_ _03832_ _03833_ _03811_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_207_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22075_ _03766_ _03767_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__nand2_1
XTAP_6749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_238_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21026_ _02790_ _02791_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__nor2_1
XFILLER_0_214_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_214_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22977_ top_inst.skew_buff_inst.row\[1\].output_reg\[7\] _04570_ VGND VGND VPWR VPWR
+ _04579_ sky130_fd_sc_hd__or2_1
XFILLER_0_214_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12730_ _05534_ _05539_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21928_ _03594_ _03642_ _03644_ _03624_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _05444_ _05445_ _05471_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__nand3_2
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21859_ _03576_ _03577_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__nand2_1
XFILLER_0_214_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14400_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[1\] _07096_ _07097_
+ VGND VGND VPWR VPWR _07098_ sky130_fd_sc_hd__and3_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15380_ _07985_ _07986_ _08023_ VGND VGND VPWR VPWR _08024_ sky130_fd_sc_hd__o21a_1
X_12592_ _05325_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_136_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24578_ clknet_leaf_142_clk _01111_ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_182_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14331_ _06995_ _07014_ _07012_ VGND VGND VPWR VPWR _07040_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23529_ clknet_leaf_139_clk net671 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17050_ _09600_ _09601_ _09595_ VGND VGND VPWR VPWR _09603_ sky130_fd_sc_hd__a21oi_1
X_14262_ _06936_ _06972_ VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_208_1124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13213_ _05989_ _05990_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16001_ _08593_ _08576_ _08609_ VGND VGND VPWR VPWR _08610_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14193_ _06857_ _06860_ _06858_ VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_221_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13144_ _05886_ _05923_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13075_ _05854_ _05855_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__nand2_1
X_17952_ _10454_ _10455_ VGND VGND VPWR VPWR _10456_ sky130_fd_sc_hd__nor2_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16903_ _09194_ _09189_ _09219_ VGND VGND VPWR VPWR _09459_ sky130_fd_sc_hd__o21a_2
X_12026_ net278 _05018_ _05029_ _05022_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__o211a_1
XFILLER_0_224_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17883_ _10338_ _10345_ _10388_ VGND VGND VPWR VPWR _10389_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_217_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19622_ _01444_ _01451_ _01452_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__nand3_1
XFILLER_0_219_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16834_ _09388_ _09389_ _09390_ VGND VGND VPWR VPWR _09392_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19553_ _06701_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__clkbuf_4
X_16765_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[5\] _09296_ _09297_
+ VGND VGND VPWR VPWR _09324_ sky130_fd_sc_hd__a21bo_1
X_13977_ _06690_ _06695_ VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18504_ _10930_ _10945_ _10965_ VGND VGND VPWR VPWR _10966_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_38_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15716_ _08324_ _08331_ VGND VGND VPWR VPWR _08332_ sky130_fd_sc_hd__xnor2_2
X_19484_ _01315_ _01316_ _01313_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__a21o_1
X_12928_ _05731_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__buf_12
X_16696_ _09247_ _09240_ _09257_ VGND VGND VPWR VPWR _09258_ sky130_fd_sc_hd__o21a_1
XFILLER_0_158_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18435_ _10897_ _10898_ VGND VGND VPWR VPWR _10899_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15647_ _05311_ VGND VGND VPWR VPWR _08265_ sky130_fd_sc_hd__buf_6
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _05664_ _05665_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__or2_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_920 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18366_ _10827_ _10829_ _10831_ VGND VGND VPWR VPWR _10832_ sky130_fd_sc_hd__o21a_1
X_15578_ _08187_ _08188_ VGND VGND VPWR VPWR _08198_ sky130_fd_sc_hd__or2b_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17317_ _09858_ _09859_ VGND VGND VPWR VPWR _09860_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14529_ _07130_ _07154_ _07155_ VGND VGND VPWR VPWR _07222_ sky130_fd_sc_hd__nand3_1
XFILLER_0_44_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18297_ _10589_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[2\] _10762_
+ _10763_ VGND VGND VPWR VPWR _10764_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17248_ _09623_ _09793_ VGND VGND VPWR VPWR _09794_ sky130_fd_sc_hd__xor2_2
XFILLER_0_153_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17179_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[15\] _09459_ _09417_
+ VGND VGND VPWR VPWR _09728_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20190_ _10030_ _11692_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__or2_2
XFILLER_0_110_842 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_243_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22900_ net771 _04522_ _04534_ _04524_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23880_ clknet_leaf_62_clk _00413_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22831_ net936 _02877_ _04495_ _03929_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22762_ _04268_ _04431_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24501_ clknet_leaf_128_clk _01034_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dfxtp_4
X_21713_ _03389_ _03392_ _03416_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__a21oi_2
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22693_ _04268_ _04349_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__nor2_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24432_ clknet_leaf_58_clk net634 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].output_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_21644_ _03210_ _03325_ _03326_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_93_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24363_ clknet_leaf_30_clk _00896_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[122\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_40 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21575_ _03305_ _03306_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__nor2_1
XANTENNA_51 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23314_ net393 _04765_ _04772_ _04769_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__o211a_1
XANTENNA_73 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20526_ _02268_ _02308_ _02309_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_84 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24294_ clknet_leaf_137_clk _00827_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_95 net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23245_ net802 _04726_ _04733_ _04730_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20457_ top_inst.grid_inst.data_path_wires\[16\]\[5\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[3\]
+ _02051_ top_inst.grid_inst.data_path_wires\[16\]\[6\] VGND VGND VPWR VPWR _02242_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23176_ net379 _04685_ _04694_ _04691_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20388_ _02174_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__clkbuf_1
XTAP_6502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22127_ _03816_ _03817_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__or2_1
XTAP_6524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22058_ _03738_ _03732_ _03750_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__nand3_1
XTAP_6579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13900_ _06632_ _06620_ VGND VGND VPWR VPWR _06633_ sky130_fd_sc_hd__or2_1
X_21009_ _02774_ _02775_ VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__or2_1
XTAP_5867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14880_ _07561_ _07563_ VGND VGND VPWR VPWR _07564_ sky130_fd_sc_hd__xor2_1
XTAP_5878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13831_ _06571_ _06556_ VGND VGND VPWR VPWR _06573_ sky130_fd_sc_hd__and2b_1
XFILLER_0_230_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16550_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[13\] _08975_ _08896_
+ VGND VGND VPWR VPWR _09126_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13762_ _06196_ _06458_ _06459_ _06421_ VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__o2bb2a_1
X_15501_ _07608_ _06634_ _08138_ _07643_ VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__o211a_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12713_ _05406_ _05522_ _05523_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__or3_1
XFILLER_0_211_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16481_ _09057_ _09058_ VGND VGND VPWR VPWR _09059_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13693_ _06436_ _06438_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18220_ _10685_ _10688_ VGND VGND VPWR VPWR _10689_ sky130_fd_sc_hd__xor2_2
XFILLER_0_35_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15432_ _08068_ _08038_ _08073_ VGND VGND VPWR VPWR _08074_ sky130_fd_sc_hd__a21oi_1
X_12644_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[3\]
+ _05287_ _05291_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__and4_1
XFILLER_0_214_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18151_ _10621_ _10622_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[1\]
+ VGND VGND VPWR VPWR _10624_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12575_ _05358_ _05388_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__xnor2_1
X_15363_ _08005_ _08006_ VGND VGND VPWR VPWR _08007_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17102_ _09611_ _09612_ VGND VGND VPWR VPWR _09654_ sky130_fd_sc_hd__or2b_1
XFILLER_0_142_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14314_ _06364_ _07023_ VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__and2_1
X_18082_ net975 _10563_ _10576_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15294_ _07901_ _07938_ VGND VGND VPWR VPWR _07940_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_230_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17033_ _09546_ _09545_ VGND VGND VPWR VPWR _09586_ sky130_fd_sc_hd__and2b_1
XFILLER_0_180_1113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14245_ _06919_ _06920_ _06917_ VGND VGND VPWR VPWR _06957_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_46_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14176_ _06856_ _06861_ _06888_ VGND VGND VPWR VPWR _06889_ sky130_fd_sc_hd__o21a_1
XFILLER_0_238_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13127_ _05903_ _05905_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18984_ _11402_ _11405_ VGND VGND VPWR VPWR _11406_ sky130_fd_sc_hd__xnor2_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _05838_ _05839_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__xor2_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ _10405_ _10406_ _10438_ VGND VGND VPWR VPWR _10440_ sky130_fd_sc_hd__and3_1
XFILLER_0_225_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12009_ net445 _05010_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__or2_1
XFILLER_0_178_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17866_ _10370_ _10369_ VGND VGND VPWR VPWR _10372_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16817_ _09371_ _09374_ VGND VGND VPWR VPWR _09375_ sky130_fd_sc_hd__xnor2_1
X_19605_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[9\] _01395_ _01396_
+ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17797_ _10303_ _10304_ VGND VGND VPWR VPWR _10305_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19536_ _01366_ _01367_ _01368_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__nand3_1
XFILLER_0_18_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16748_ _09211_ _09187_ _09306_ _09307_ VGND VGND VPWR VPWR _09308_ sky130_fd_sc_hd__and4_1
XFILLER_0_117_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19467_ _11678_ _11705_ _11708_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__and3_1
XFILLER_0_220_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16679_ _09240_ _09241_ VGND VGND VPWR VPWR _09242_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18418_ _10867_ _10869_ VGND VGND VPWR VPWR _10882_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19398_ _01213_ _01215_ _01232_ _01233_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18349_ _10761_ _10773_ VGND VGND VPWR VPWR _10815_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21360_ _03088_ _03096_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__xor2_2
XFILLER_0_71_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20311_ _02068_ _02094_ _02096_ _02070_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_163_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold800 top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[6\] VGND VGND
+ VPWR VPWR net982 sky130_fd_sc_hd__dlygate4sd3_1
X_21291_ _03028_ _03029_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold811 top_inst.axis_out_inst.out_buff_data\[99\] VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23030_ net616 _04603_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__or2_1
Xhold822 top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[1\] VGND VGND
+ VPWR VPWR net1004 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold833 top_inst.axis_in_inst.inbuf_bus\[23\] VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__dlygate4sd3_1
X_20242_ _02032_ _02033_ _06178_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__o21ai_1
Xhold844 top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[1\] VGND VGND
+ VPWR VPWR net1026 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold855 top_inst.axis_in_inst.inbuf_bus\[22\] VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold866 top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[3\] VGND VGND
+ VPWR VPWR net1048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold877 top_inst.axis_out_inst.out_buff_data\[61\] VGND VGND VPWR VPWR net1059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold888 top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[4\] VGND VGND
+ VPWR VPWR net1070 sky130_fd_sc_hd__dlygate4sd3_1
X_20173_ _01964_ _01969_ _01982_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_228_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold899 top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[4\] VGND VGND
+ VPWR VPWR net1081 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23932_ clknet_leaf_91_clk _00465_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23863_ clknet_leaf_68_clk _00396_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_211_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22814_ _04411_ _04430_ _04268_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23794_ clknet_leaf_69_clk _00327_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22745_ _04388_ _04392_ _04414_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__nand3_1
XFILLER_0_149_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22676_ _04137_ _04331_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24415_ clknet_leaf_56_clk _00948_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21627_ _03351_ _03355_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_192_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12360_ net300 _05209_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__or2_1
X_24346_ clknet_leaf_24_clk _00879_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[105\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21558_ _03253_ _03289_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_209_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_1299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20509_ _02287_ _02244_ _02290_ _02291_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__or4_2
XFILLER_0_121_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12291_ net466 _05169_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__or2_1
X_24277_ clknet_leaf_11_clk _00810_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[17\]\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_106_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21489_ _03207_ _03222_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__xor2_2
XFILLER_0_50_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14030_ _06745_ _06746_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23228_ net651 _04713_ _04723_ _04717_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__o211a_1
XFILLER_0_240_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23159_ net76 _04672_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15981_ _08588_ _08590_ _06734_ VGND VGND VPWR VPWR _08591_ sky130_fd_sc_hd__a21oi_1
XTAP_5631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17720_ _10229_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14932_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[31\] _07576_ VGND
+ VGND VPWR VPWR _07605_ sky130_fd_sc_hd__and2_1
XTAP_5664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ _10037_ top_inst.grid_inst.data_path_wires\[11\]\[5\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _10162_ sky130_fd_sc_hd__nand4_1
XFILLER_0_215_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14863_ _07514_ _07547_ VGND VGND VPWR VPWR _07548_ sky130_fd_sc_hd__or2_1
XTAP_4963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16602_ _09055_ _09153_ _09152_ VGND VGND VPWR VPWR _09176_ sky130_fd_sc_hd__o21a_1
XTAP_4996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13814_ _06537_ _06541_ _06535_ VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__o21a_1
X_17582_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[2\] _10073_ _10074_
+ VGND VGND VPWR VPWR _10096_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_202_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14794_ _07444_ _07479_ VGND VGND VPWR VPWR _07481_ sky130_fd_sc_hd__or2_1
XFILLER_0_212_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19321_ _11684_ _11679_ _11677_ _11682_ VGND VGND VPWR VPWR _11716_ sky130_fd_sc_hd__nand4_1
XFILLER_0_97_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16533_ _09108_ _09109_ VGND VGND VPWR VPWR _09110_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13745_ _06196_ _06212_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19252_ _11514_ _11648_ _11665_ VGND VGND VPWR VPWR _11666_ sky130_fd_sc_hd__o21a_1
X_16464_ _08697_ _08676_ _09041_ VGND VGND VPWR VPWR _09042_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13676_ _06420_ _06421_ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__xor2_1
XFILLER_0_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18203_ _10608_ _10645_ _10672_ VGND VGND VPWR VPWR _10673_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_26_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15415_ _08055_ _08057_ VGND VGND VPWR VPWR _08058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19183_ _11164_ _11598_ _11559_ _11599_ VGND VGND VPWR VPWR _11600_ sky130_fd_sc_hd__a22oi_2
X_12627_ _04867_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__buf_8
XFILLER_0_109_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16395_ _08897_ VGND VGND VPWR VPWR _08975_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18134_ _10610_ _10057_ VGND VGND VPWR VPWR _10611_ sky130_fd_sc_hd__or2_1
X_15346_ _07624_ _07637_ VGND VGND VPWR VPWR _07990_ sky130_fd_sc_hd__nand2_2
X_12558_ _05350_ _05371_ _05315_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18065_ _10546_ _10552_ _10554_ VGND VGND VPWR VPWR _10565_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15277_ _07921_ _07922_ VGND VGND VPWR VPWR _07923_ sky130_fd_sc_hd__nor2_1
X_12489_ _05304_ _05276_ _05307_ _05308_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold107 _00289_ VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold118 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[31\] VGND
+ VGND VPWR VPWR net300 sky130_fd_sc_hd__dlygate4sd3_1
X_17016_ _09567_ _09568_ _09521_ _09543_ VGND VGND VPWR VPWR _09570_ sky130_fd_sc_hd__o211ai_2
Xhold129 top_inst.deskew_buff_inst.col_input\[16\] VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__dlygate4sd3_1
X_14228_ _06938_ _06901_ _06939_ VGND VGND VPWR VPWR _06940_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14159_ _06822_ _06820_ VGND VGND VPWR VPWR _06873_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18967_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[9\] _11340_ VGND
+ VGND VPWR VPWR _11389_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_226_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17918_ _10419_ _10421_ _10422_ VGND VGND VPWR VPWR _10423_ sky130_fd_sc_hd__nor3_1
X_18898_ _11307_ _11321_ VGND VGND VPWR VPWR _11322_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_240_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17849_ _10354_ _10355_ VGND VGND VPWR VPWR _10356_ sky130_fd_sc_hd__and2_1
XFILLER_0_234_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20860_ _02589_ _02611_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19519_ _11683_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[0\] _11708_
+ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20791_ _02546_ _02542_ _02565_ _01984_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22530_ _04188_ _04210_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__or2b_1
XFILLER_0_232_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22461_ _04134_ _04143_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_228_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21412_ _03145_ _03147_ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__xnor2_2
X_24200_ clknet_leaf_117_clk _00733_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22392_ _04025_ _04033_ _04076_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24131_ clknet_leaf_119_clk _00664_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_115_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21343_ _03079_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24062_ clknet_leaf_84_clk _00595_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold630 top_inst.deskew_buff_inst.col_input\[5\] VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__dlygate4sd3_1
X_21274_ _03011_ _03012_ _02871_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[2\]
+ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_163_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold641 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[30\] VGND
+ VGND VPWR VPWR net823 sky130_fd_sc_hd__dlygate4sd3_1
X_23013_ top_inst.skew_buff_inst.row\[0\].output_reg\[7\] _04596_ VGND VGND VPWR VPWR
+ _04599_ sky130_fd_sc_hd__or2_1
Xhold652 top_inst.deskew_buff_inst.col_input\[110\] VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold663 top_inst.axis_out_inst.out_buff_data\[38\] VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__dlygate4sd3_1
X_20225_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _02020_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_198_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold674 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[13\] VGND
+ VGND VPWR VPWR net856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold685 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[1\] VGND VGND
+ VPWR VPWR net867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold696 top_inst.deskew_buff_inst.col_input\[83\] VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_239_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20156_ _01924_ _01927_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20087_ _01899_ _01900_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__nand2_1
XTAP_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23915_ clknet_leaf_33_clk _00448_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ net803 _04930_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__or2_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23846_ clknet_leaf_95_clk _00379_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11791_ net866 _04885_ _04895_ _04889_ VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__o211a_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23777_ clknet_leaf_64_clk _00310_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20989_ _02730_ _02756_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13530_ _06244_ _06248_ _06247_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__o21ba_1
X_22728_ _04349_ _04396_ _04399_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13461_ _06198_ _06204_ _06216_ _06207_ VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22659_ _04315_ _04328_ _04333_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15200_ _07788_ _07790_ _07846_ VGND VGND VPWR VPWR _07848_ sky130_fd_sc_hd__and3_1
X_12412_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[21\] _05248_
+ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16180_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[8\]\[2\]
+ top_inst.grid_inst.data_path_wires\[8\]\[1\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[4\]
+ VGND VGND VPWR VPWR _08765_ sky130_fd_sc_hd__a22o_1
X_13392_ _06136_ _06141_ _06163_ _05405_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_106_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15131_ _07747_ _07752_ VGND VGND VPWR VPWR _07780_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12343_ net321 _05209_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__or2_1
X_24329_ clknet_leaf_6_clk _00862_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15062_ top_inst.grid_inst.data_path_wires\[6\]\[2\] top_inst.grid_inst.data_path_wires\[6\]\[1\]
+ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _07713_ sky130_fd_sc_hd__nand4_4
X_12274_ net976 _05164_ _05171_ _05168_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14013_ _06704_ _06729_ _05399_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19870_ _01678_ _01693_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18821_ _11230_ _11246_ VGND VGND VPWR VPWR _11247_ sky130_fd_sc_hd__xor2_2
XTAP_6140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18752_ _11179_ _11180_ VGND VGND VPWR VPWR _11181_ sky130_fd_sc_hd__nand2_1
XTAP_5450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15964_ _08572_ _08573_ VGND VGND VPWR VPWR _08574_ sky130_fd_sc_hd__nor2_1
XTAP_6195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17703_ _10211_ _10212_ VGND VGND VPWR VPWR _10213_ sky130_fd_sc_hd__xnor2_1
X_14915_ net229 _07596_ _07594_ VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__o21a_1
XTAP_5483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18683_ top_inst.grid_inst.data_path_wires\[13\]\[0\] VGND VGND VPWR VPWR _11130_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_234_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15895_ _08453_ _08456_ _08506_ VGND VGND VPWR VPWR _08507_ sky130_fd_sc_hd__a21bo_1
XTAP_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_231_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_1175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17634_ _10143_ _10145_ VGND VGND VPWR VPWR _10146_ sky130_fd_sc_hd__xnor2_2
X_14846_ _07415_ VGND VGND VPWR VPWR _07531_ sky130_fd_sc_hd__inv_2
XTAP_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17565_ _10072_ _10078_ VGND VGND VPWR VPWR _10080_ sky130_fd_sc_hd__nand2_1
X_14777_ _07459_ _07463_ VGND VGND VPWR VPWR _07464_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11989_ net722 _05004_ _05007_ _05008_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19304_ _05755_ _11700_ _11702_ _11641_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16516_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[12\] _08975_ _08896_
+ VGND VGND VPWR VPWR _09093_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13728_ _06470_ _06472_ VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__xor2_1
X_17496_ top_inst.grid_inst.data_path_wires\[11\]\[2\] VGND VGND VPWR VPWR _10027_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19235_ _11647_ _11649_ VGND VGND VPWR VPWR _11650_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16447_ _09020_ _09025_ VGND VGND VPWR VPWR _09026_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13659_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[8\] _06242_ _06403_
+ _06405_ VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19166_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[13\] _10364_ _11582_
+ _11583_ _11228_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16378_ _08926_ _08925_ VGND VGND VPWR VPWR _08958_ sky130_fd_sc_hd__or2b_1
XFILLER_0_60_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18117_ _10577_ _10046_ _10598_ _10594_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15329_ _07972_ _07973_ VGND VGND VPWR VPWR _07974_ sky130_fd_sc_hd__xnor2_2
X_19097_ _11514_ _11515_ VGND VGND VPWR VPWR _11516_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18048_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[16\] _10367_ VGND
+ VGND VPWR VPWR _10549_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_223_1035 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_240_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20010_ _01801_ _01804_ _01803_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19999_ _01798_ _01816_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__nor2_1
XFILLER_0_193_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21961_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[31\] _03669_ VGND
+ VGND VPWR VPWR _03675_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23700_ clknet_leaf_125_clk _00233_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20912_ top_inst.deskew_buff_inst.col_input\[54\] _11723_ _02664_ _02682_ VGND VGND
+ VPWR VPWR _02683_ sky130_fd_sc_hd__a22o_1
X_21892_ _03610_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23631_ clknet_leaf_102_clk net507 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_20843_ _02463_ _02601_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_230_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23562_ clknet_leaf_100_clk net815 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_20774_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[17\] _02467_ VGND
+ VGND VPWR VPWR _02550_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22513_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[15\] _03937_ _03938_
+ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23493_ clknet_leaf_142_clk _00026_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[83\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22444_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[13\] _03937_ _03938_
+ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22375_ _03950_ _04023_ _03983_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24114_ clknet_leaf_16_clk _00647_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21326_ _03024_ _03063_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__xor2_1
XFILLER_0_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24045_ clknet_leaf_42_clk _00578_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold460 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[1\] VGND
+ VGND VPWR VPWR net642 sky130_fd_sc_hd__dlygate4sd3_1
X_21257_ _02972_ _02978_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__or2b_1
Xhold471 top_inst.valid_pipe\[4\] VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold482 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[30\] VGND
+ VGND VPWR VPWR net664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 _00907_ VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20208_ _01987_ _11163_ _02008_ _02006_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21188_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[3\] _02928_ _02929_
+ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__and3_1
XFILLER_0_244_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20139_ _01934_ _01937_ _01936_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12961_ _05755_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__clkbuf_4
XTAP_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14700_ _07371_ _07387_ _07388_ VGND VGND VPWR VPWR _07389_ sky130_fd_sc_hd__nand3_1
XFILLER_0_169_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _04911_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__clkbuf_4
XTAP_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15680_ _08295_ _08293_ _08294_ VGND VGND VPWR VPWR _08297_ sky130_fd_sc_hd__and3_1
XTAP_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _05352_ _05697_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _07070_ _07086_ _07288_ _07287_ VGND VGND VPWR VPWR _07321_ sky130_fd_sc_hd__a31o_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23829_ clknet_leaf_93_clk _00362_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_11843_ _04911_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__clkbuf_4
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17350_ _09882_ _09889_ _09887_ _09890_ VGND VGND VPWR VPWR _09891_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_71_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _07251_ _07252_ _07234_ VGND VGND VPWR VPWR _07254_ sky130_fd_sc_hd__a21o_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ net377 _04877_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _08880_ _08882_ VGND VGND VPWR VPWR _08883_ sky130_fd_sc_hd__xnor2_2
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _06250_ _06255_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__and2_1
X_17281_ _09767_ _09823_ _09825_ _09800_ VGND VGND VPWR VPWR _09826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14493_ _07130_ _07155_ _07186_ VGND VGND VPWR VPWR _07187_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19020_ _11400_ _11440_ VGND VGND VPWR VPWR _11441_ sky130_fd_sc_hd__xor2_1
X_16232_ _08806_ _08814_ VGND VGND VPWR VPWR _08816_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13444_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _06205_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_222_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16163_ _08747_ _08748_ VGND VGND VPWR VPWR _08749_ sky130_fd_sc_hd__xnor2_2
X_13375_ _06085_ _06116_ _06117_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_140_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15114_ _07754_ _07763_ VGND VGND VPWR VPWR _07764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12326_ net480 _05196_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__or2_1
X_16094_ _08667_ _08681_ _08689_ _08666_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19922_ _01738_ _01742_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__xor2_4
X_15045_ top_inst.grid_inst.data_path_wires\[6\]\[0\] _07635_ _07633_ top_inst.grid_inst.data_path_wires\[6\]\[1\]
+ VGND VGND VPWR VPWR _07697_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12257_ net435 _05151_ _05161_ _05155_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12188_ net836 _05110_ _05121_ _05114_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__o211a_1
X_19853_ _11177_ _01676_ _01677_ _11714_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__o211a_1
X_18804_ _11216_ _11221_ VGND VGND VPWR VPWR _11230_ sky130_fd_sc_hd__and2b_1
XFILLER_0_194_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16996_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[4\] _09203_ _09218_
+ VGND VGND VPWR VPWR _09550_ sky130_fd_sc_hd__o21ai_2
X_19784_ _01486_ _01487_ _01606_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_207_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18735_ _11147_ _11163_ _11166_ _11160_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__o211a_1
X_15947_ _08522_ _08523_ VGND VGND VPWR VPWR _08557_ sky130_fd_sc_hd__nand2_1
XTAP_5280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18666_ _11121_ _11122_ VGND VGND VPWR VPWR _11123_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ _08438_ _08440_ _08437_ VGND VGND VPWR VPWR _08490_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_91_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14829_ _07485_ _07475_ _07513_ VGND VGND VPWR VPWR _07515_ sky130_fd_sc_hd__or3_1
XFILLER_0_203_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17617_ top_inst.grid_inst.data_path_wires\[11\]\[2\] top_inst.grid_inst.data_path_wires\[11\]\[1\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[4\] VGND VGND VPWR VPWR
+ _10129_ sky130_fd_sc_hd__and3_1
XFILLER_0_231_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18597_ _10933_ _11056_ VGND VGND VPWR VPWR _11057_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17548_ top_inst.grid_inst.data_path_wires\[11\]\[0\] _10044_ _10042_ _10025_ VGND
+ VGND VPWR VPWR _10064_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_1311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17479_ _10013_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19218_ _11587_ _11609_ _11607_ VGND VGND VPWR VPWR _11634_ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20490_ _02231_ _02233_ VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19149_ _11479_ _11565_ VGND VGND VPWR VPWR _11567_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22160_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[6\] _03814_ _03815_
+ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21111_ _06619_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__buf_2
XFILLER_0_160_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22091_ _03781_ _03782_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21042_ _02710_ _02712_ _02714_ _02806_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_227_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1062 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22993_ net583 _04575_ _04587_ _04577_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21944_ _02706_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21875_ _03563_ _03566_ _03589_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_221_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23614_ clknet_leaf_105_clk _00147_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_20826_ _02598_ _02599_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__nor2_1
XFILLER_0_194_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24594_ clknet_leaf_22_clk _01127_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_33_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23545_ clknet_leaf_129_clk _00078_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_143_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_143_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20757_ _02532_ _02533_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23476_ clknet_leaf_136_clk _00009_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20688_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[7\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[4\]
+ _02003_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__mux2_4
XFILLER_0_123_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22427_ _04108_ _04110_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13160_ _05937_ _05938_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22358_ _03977_ _04002_ _04043_ VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_131_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12111_ net254 _05071_ _05078_ _05075_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__o211a_1
X_13091_ _05863_ _05871_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21309_ _03045_ _03046_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22289_ _03936_ _03967_ _03975_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_1375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12042_ net510 _05036_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__or2_1
X_24028_ clknet_leaf_48_clk _00561_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold290 _00005_ VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16850_ _08831_ _09407_ VGND VGND VPWR VPWR _09408_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15801_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[8\] _08374_ _08373_
+ VGND VGND VPWR VPWR _08415_ sky130_fd_sc_hd__a21o_1
XFILLER_0_232_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16781_ _09335_ _09336_ _09339_ VGND VGND VPWR VPWR _09340_ sky130_fd_sc_hd__nand3_1
XFILLER_0_189_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13993_ _06626_ _06643_ _06709_ _06710_ VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_244_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18520_ _10934_ _10936_ VGND VGND VPWR VPWR _10982_ sky130_fd_sc_hd__nor2_1
XFILLER_0_232_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15732_ _08347_ VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__clkbuf_1
X_12944_ top_inst.grid_inst.data_path_wires\[1\]\[3\] VGND VGND VPWR VPWR _05744_
+ sky130_fd_sc_hd__buf_4
XFILLER_0_77_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18451_ _10874_ _10913_ VGND VGND VPWR VPWR _10915_ sky130_fd_sc_hd__or2_1
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ _08163_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[2\] _08277_
+ _08278_ VGND VGND VPWR VPWR _08280_ sky130_fd_sc_hd__nand4_2
X_12875_ _05608_ _05679_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__or2_1
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17402_ _09913_ _09934_ _09939_ VGND VGND VPWR VPWR _09941_ sky130_fd_sc_hd__nand3_1
XFILLER_0_158_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _07275_ _07304_ VGND VGND VPWR VPWR _07305_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _10808_ _10806_ VGND VGND VPWR VPWR _10847_ sky130_fd_sc_hd__or2b_1
X_11826_ _04874_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__clkbuf_4
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _08195_ _08212_ _08213_ VGND VGND VPWR VPWR _08214_ sky130_fd_sc_hd__or3_1
XFILLER_0_200_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17333_ _09624_ _09873_ VGND VGND VPWR VPWR _09875_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _07079_ _07073_ _07077_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _07237_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_173_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_134_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_134_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11757_ _04863_ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_166_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17264_ _09726_ _09795_ VGND VGND VPWR VPWR _09809_ sky130_fd_sc_hd__nor2_1
X_14476_ _07167_ _07168_ _07162_ VGND VGND VPWR VPWR _07170_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19003_ _11382_ _11423_ _09292_ VGND VGND VPWR VPWR _11425_ sky130_fd_sc_hd__a21o_1
X_16215_ _08797_ _08798_ VGND VGND VPWR VPWR _08799_ sky130_fd_sc_hd__nand2_1
X_13427_ top_inst.grid_inst.data_path_wires\[2\]\[5\] VGND VGND VPWR VPWR _06193_
+ sky130_fd_sc_hd__buf_4
X_17195_ _09721_ _09743_ VGND VGND VPWR VPWR _09744_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16146_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[2\] _08711_ _08712_
+ VGND VGND VPWR VPWR _08733_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13358_ _06130_ _06131_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_224_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12309_ _05177_ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__buf_2
X_16077_ _08676_ VGND VGND VPWR VPWR _08677_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13289_ _05945_ _06064_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_922 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19905_ _01611_ _01701_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__nor2_1
X_15028_ _07668_ _07662_ _07680_ VGND VGND VPWR VPWR _07681_ sky130_fd_sc_hd__a21o_1
XFILLER_0_220_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19836_ _01528_ _01659_ _01660_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_78_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19767_ _01560_ _01554_ _01590_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__a21oi_1
X_16979_ _09409_ _09449_ _09492_ _09533_ VGND VGND VPWR VPWR _09534_ sky130_fd_sc_hd__o31ai_1
Xinput3 input_tdata[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_194_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18718_ _11154_ _11150_ VGND VGND VPWR VPWR _11155_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_1370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19698_ _01402_ _01485_ _01484_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_231_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_235_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18649_ _11079_ _11082_ _11106_ VGND VGND VPWR VPWR _11107_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_231_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21660_ _03387_ _03388_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__or2_2
XFILLER_0_176_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20611_ _02354_ _02377_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_125_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_125_clk
+ sky130_fd_sc_hd__clkbuf_16
X_21591_ _03210_ _03294_ _03321_ VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_149_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23330_ _04690_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__buf_4
XFILLER_0_74_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20542_ _01997_ _02188_ _02324_ _02186_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1027 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23261_ _04690_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__buf_4
X_20473_ _02255_ _02256_ _02224_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22212_ _03693_ _03703_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23192_ _04690_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22143_ _03811_ _03832_ _03833_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1094 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22074_ _03705_ top_inst.grid_inst.data_path_wires\[18\]\[1\] top_inst.grid_inst.data_path_wires\[18\]\[0\]
+ _03707_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__a22o_1
XTAP_6739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21025_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[25\] _02559_ _02789_
+ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_242_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22976_ net637 _04575_ _04578_ _04577_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21927_ _03611_ _03607_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__nand2_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_214_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _05444_ _05445_ _05471_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__a21o_2
XFILLER_0_84_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21858_ _03576_ _03577_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20809_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[16\] _02559_ _02553_
+ _02551_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12591_ net982 _05403_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__nand2_1
X_24577_ clknet_leaf_140_clk _01110_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_116_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21789_ _03478_ _03511_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__nand2_1
XFILLER_0_203_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14330_ _06995_ _07038_ VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_943 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23528_ clknet_leaf_139_clk _00061_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14261_ _06970_ _06971_ VGND VGND VPWR VPWR _06972_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23459_ top_inst.axis_out_inst.out_buff_data\[117\] _04864_ VGND VGND VPWR VPWR _04852_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_208_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16000_ _08602_ _08608_ VGND VGND VPWR VPWR _08609_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_208_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13212_ _05945_ _05988_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14192_ _06903_ _06904_ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_979 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13143_ _05887_ _05920_ _05921_ _05922_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _05738_ top_inst.grid_inst.data_path_wires\[1\]\[0\] _05770_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[5\]
+ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__nand4_2
X_17951_ _10413_ _10453_ VGND VGND VPWR VPWR _10455_ sky130_fd_sc_hd__and2_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16902_ _09422_ _09439_ _09440_ VGND VGND VPWR VPWR _09458_ sky130_fd_sc_hd__nand3_1
X_12025_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[15\] _05023_
+ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__or2_1
X_17882_ _10344_ _10343_ VGND VGND VPWR VPWR _10388_ sky130_fd_sc_hd__or2b_1
XFILLER_0_79_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19621_ _01448_ _01449_ _01450_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__a21o_1
XFILLER_0_217_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16833_ _09388_ _09389_ _09390_ VGND VGND VPWR VPWR _09391_ sky130_fd_sc_hd__and3_1
XFILLER_0_232_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16764_ _09323_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__clkbuf_1
X_19552_ _01345_ net210 VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__xor2_2
X_13976_ _06691_ _06694_ VGND VGND VPWR VPWR _06695_ sky130_fd_sc_hd__xor2_1
XFILLER_0_232_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15715_ _08329_ _08330_ VGND VGND VPWR VPWR _08331_ sky130_fd_sc_hd__nor2_1
X_18503_ _10942_ _10944_ VGND VGND VPWR VPWR _10965_ sky130_fd_sc_hd__and2b_1
XFILLER_0_232_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12927_ _05730_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__buf_6
X_16695_ _09253_ _09256_ VGND VGND VPWR VPWR _09257_ sky130_fd_sc_hd__xnor2_1
X_19483_ _01313_ _01315_ _01316_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18434_ top_inst.grid_inst.data_path_wires\[12\]\[4\] _10612_ _10857_ top_inst.grid_inst.data_path_wires\[12\]\[3\]
+ VGND VGND VPWR VPWR _10898_ sky130_fd_sc_hd__o2bb2a_1
X_15646_ _08237_ _08263_ VGND VGND VPWR VPWR _08264_ sky130_fd_sc_hd__nand2_1
X_12858_ _05636_ _05624_ _05663_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18365_ _05310_ VGND VGND VPWR VPWR _10831_ sky130_fd_sc_hd__buf_8
XFILLER_0_16_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11809_ top_inst.axis_out_inst.out_buff_data\[82\] _04903_ VGND VGND VPWR VPWR _04906_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_173_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15577_ _04869_ VGND VGND VPWR VPWR _08197_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_107_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_200_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12789_ _05296_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _09833_ _09841_ _09856_ _09816_ VGND VGND VPWR VPWR _09859_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14528_ _07219_ _07220_ VGND VGND VPWR VPWR _07221_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18296_ _10606_ _10585_ _10608_ _10604_ VGND VGND VPWR VPWR _10763_ sky130_fd_sc_hd__nand4_2
XFILLER_0_84_896 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17247_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[19\] _09631_ VGND
+ VGND VPWR VPWR _09793_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14459_ net1125 _07152_ _07153_ VGND VGND VPWR VPWR _07154_ sky130_fd_sc_hd__or3b_2
XFILLER_0_142_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17178_ _09726_ _09706_ _09677_ VGND VGND VPWR VPWR _09727_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_12_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16129_ _08710_ _08716_ VGND VGND VPWR VPWR _08717_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19819_ _01628_ _01644_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22830_ top_inst.skew_buff_inst.row\[3\].output_reg\[0\] _03691_ VGND VGND VPWR VPWR
+ _04495_ sky130_fd_sc_hd__or2_1
XFILLER_0_211_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22761_ _04410_ _04430_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_17_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24500_ clknet_leaf_126_clk _01033_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_220_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21712_ _03394_ _03417_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__or2b_1
XFILLER_0_17_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22692_ _04351_ _04344_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24431_ clknet_leaf_58_clk net638 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].output_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21643_ _03352_ _03354_ _03371_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24362_ clknet_leaf_30_clk _00895_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[121\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_30 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21574_ _03302_ _03304_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_41 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_52 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_244_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_63 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23313_ net148 _04766_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20525_ _02268_ _02308_ _07576_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__a21oi_1
XANTENNA_74 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24293_ clknet_leaf_120_clk _00826_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_85 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23244_ net115 _04727_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__or2_1
X_20456_ _02003_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[1\] VGND
+ VGND VPWR VPWR _02241_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1058 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23175_ net82 _04687_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__or2_1
X_20387_ _02135_ _02173_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__and2_1
XFILLER_0_219_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22126_ _03814_ _03815_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[6\]
+ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22057_ _03738_ _03732_ _03750_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__a21o_1
XTAP_5835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21008_ _02749_ _02764_ _02773_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__and3_1
XTAP_5868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13830_ _06556_ _06571_ VGND VGND VPWR VPWR _06572_ sky130_fd_sc_hd__and2b_1
XFILLER_0_216_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_230_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_1274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13761_ _06503_ _06504_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__nor2_1
X_22959_ net404 _04562_ _04568_ _04564_ VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15500_ _08137_ _06620_ VGND VGND VPWR VPWR _08138_ sky130_fd_sc_hd__or2_1
X_12712_ _05520_ _05521_ _05476_ _05479_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16480_ _09055_ _09056_ VGND VGND VPWR VPWR _09058_ sky130_fd_sc_hd__and2_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13692_ _06390_ _06437_ _06387_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__o21a_1
XFILLER_0_214_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15431_ _07956_ _08072_ VGND VGND VPWR VPWR _08073_ sky130_fd_sc_hd__xor2_1
XFILLER_0_210_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12643_ _05293_ _05287_ _05292_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_182_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24629_ clknet_leaf_22_clk _01162_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[105\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_1436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18150_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[1\] _10621_ _10622_
+ VGND VGND VPWR VPWR _10623_ sky130_fd_sc_hd__nand3_1
XFILLER_0_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15362_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[12\] _07845_ VGND
+ VGND VPWR VPWR _08006_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12574_ _05384_ _05387_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_1211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17101_ _09627_ _09652_ VGND VGND VPWR VPWR _09653_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_136_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14313_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[13\] _07022_ _06701_
+ VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18081_ net961 _10563_ _10576_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__o21a_1
XFILLER_0_230_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15293_ _07901_ _07938_ VGND VGND VPWR VPWR _07939_ sky130_fd_sc_hd__and2_1
X_17032_ _09542_ _09570_ _09569_ VGND VGND VPWR VPWR _09585_ sky130_fd_sc_hd__a21bo_1
X_14244_ _06953_ _06955_ VGND VGND VPWR VPWR _06956_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_230_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_1125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14175_ _06855_ _06854_ VGND VGND VPWR VPWR _06888_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13126_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[7\] _05903_ _05905_
+ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ _11403_ _11404_ VGND VGND VPWR VPWR _11405_ sky130_fd_sc_hd__nor2_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _05803_ _05807_ _05806_ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__o21ba_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _10405_ _10406_ _10438_ VGND VGND VPWR VPWR _10439_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12008_ net745 _05018_ _05019_ _05008_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_1140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17865_ _10369_ _10370_ VGND VGND VPWR VPWR _10371_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_233_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19604_ _01401_ _01418_ _01419_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__nand3_1
X_16816_ _09372_ _09373_ VGND VGND VPWR VPWR _09374_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17796_ _10029_ _10054_ _10248_ _10247_ VGND VGND VPWR VPWR _10304_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_233_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19535_ _01313_ _01316_ _01315_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__a21bo_1
X_16747_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[2\] _09202_ _09304_
+ _09305_ VGND VGND VPWR VPWR _09307_ sky130_fd_sc_hd__a22o_1
X_13959_ _06667_ _06678_ VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_242_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16678_ _09232_ _09239_ VGND VGND VPWR VPWR _09241_ sky130_fd_sc_hd__and2_1
X_19466_ _01271_ _01272_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_158_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18417_ _10836_ _10876_ _10880_ _10835_ VGND VGND VPWR VPWR _10881_ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15629_ _08245_ _08246_ VGND VGND VPWR VPWR _08247_ sky130_fd_sc_hd__and2_1
X_19397_ _01230_ _01231_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[5\]
+ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18348_ _10796_ _10813_ VGND VGND VPWR VPWR _10814_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_228_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18279_ _10745_ _10746_ VGND VGND VPWR VPWR _10747_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20310_ _02075_ _02098_ _04870_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21290_ _02936_ _02958_ _02984_ _02988_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__o31a_1
XFILLER_0_86_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold801 top_inst.axis_in_inst.inbuf_bus\[1\] VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold812 top_inst.axis_in_inst.inbuf_bus\[18\] VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold823 top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[2\] VGND VGND
+ VPWR VPWR net1005 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20241_ _02024_ _02030_ _02031_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold834 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[9\] VGND VGND
+ VPWR VPWR net1016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold845 top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[1\] VGND VGND
+ VPWR VPWR net1027 sky130_fd_sc_hd__buf_1
XFILLER_0_25_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold856 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[11\] VGND VGND
+ VPWR VPWR net1038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[13\] VGND VGND
+ VPWR VPWR net1049 sky130_fd_sc_hd__dlygate4sd3_1
X_20172_ _01974_ _01981_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__xnor2_2
Xhold878 top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[1\] VGND VGND
+ VPWR VPWR net1060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold889 top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[4\] VGND VGND
+ VPWR VPWR net1071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_243_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23931_ clknet_leaf_75_clk _00464_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23862_ clknet_leaf_68_clk _00395_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22813_ _04479_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23793_ clknet_leaf_71_clk _00326_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_135_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22744_ _04388_ _04392_ _04414_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__a21o_1
XFILLER_0_211_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_211_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22675_ _04330_ _04348_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_149_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24414_ clknet_leaf_56_clk _00947_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21626_ _03351_ _03355_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24345_ clknet_leaf_24_clk _00878_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[104\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21557_ _03287_ _03288_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_181_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20508_ _02287_ _02244_ _02290_ _02291_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__o22ai_2
X_12290_ net589 _05178_ _05180_ _05168_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__o211a_1
X_24276_ clknet_leaf_11_clk _00809_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[17\]\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_181_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21488_ _03219_ _03221_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_209_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23227_ net107 _04714_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20439_ _01993_ _02016_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[6\]
+ _02184_ _02223_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__a41o_1
XFILLER_0_120_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23158_ net774 _04671_ _04682_ _04675_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__o211a_1
XTAP_6311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22109_ _03798_ _03800_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__xnor2_1
XTAP_6344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15980_ _08549_ _08551_ _08589_ VGND VGND VPWR VPWR _08590_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_101_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23089_ _04550_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_235_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14931_ _07593_ _07604_ _07594_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__o21a_1
XTAP_5643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14862_ _07520_ _07546_ VGND VGND VPWR VPWR _07547_ sky130_fd_sc_hd__xor2_1
XTAP_5698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17650_ top_inst.grid_inst.data_path_wires\[11\]\[5\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[0\] _10037_ VGND VGND
+ VPWR VPWR _10161_ sky130_fd_sc_hd__a22o_1
XTAP_4964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_215_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16601_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[15\] _08975_ _08896_
+ VGND VGND VPWR VPWR _09175_ sky130_fd_sc_hd__a21o_1
XTAP_4986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13813_ _06539_ VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__inv_2
XFILLER_0_230_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17581_ _10093_ _10094_ VGND VGND VPWR VPWR _10095_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14793_ _07444_ _07479_ VGND VGND VPWR VPWR _07480_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16532_ _09105_ _09107_ VGND VGND VPWR VPWR _09109_ sky130_fd_sc_hd__or2_1
X_19320_ _11684_ _11677_ _11682_ _11679_ VGND VGND VPWR VPWR _11715_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13744_ _06486_ _06487_ VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19251_ _11514_ _11648_ _11647_ VGND VGND VPWR VPWR _11665_ sky130_fd_sc_hd__a21o_1
X_16463_ _08876_ _08673_ VGND VGND VPWR VPWR _09041_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13675_ _06198_ _06205_ VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__nand2_2
XFILLER_0_195_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15414_ _08011_ _08012_ _08056_ VGND VGND VPWR VPWR _08057_ sky130_fd_sc_hd__a21bo_1
X_18202_ top_inst.grid_inst.data_path_wires\[12\]\[0\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[12\]\[1\]
+ VGND VGND VPWR VPWR _10672_ sky130_fd_sc_hd__a22o_1
XPHY_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12626_ _05406_ _05437_ _05438_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__or3_1
X_19182_ _11598_ _11561_ VGND VGND VPWR VPWR _11599_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16394_ _08972_ _08973_ VGND VGND VPWR VPWR _08974_ sky130_fd_sc_hd__nor2_1
XPHY_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18133_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _10610_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_183_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15345_ _07963_ _07962_ VGND VGND VPWR VPWR _07989_ sky130_fd_sc_hd__or2b_1
XFILLER_0_124_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12557_ _05350_ _05371_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_721 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18064_ _10556_ _10558_ VGND VGND VPWR VPWR _10564_ sky130_fd_sc_hd__nor2_1
X_15276_ _07920_ _07908_ VGND VGND VPWR VPWR _07922_ sky130_fd_sc_hd__and2b_1
XFILLER_0_124_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12488_ _05260_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__buf_4
Xhold108 top_inst.deskew_buff_inst.col_input\[103\] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dlygate4sd3_1
X_17015_ _09521_ _09543_ _09567_ _09568_ VGND VGND VPWR VPWR _09569_ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14227_ _06896_ _06895_ VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__and2b_1
Xhold119 _00294_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14158_ _06866_ _06871_ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13109_ top_inst.grid_inst.data_path_wires\[1\]\[1\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14089_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[7\] _05634_ _06803_
+ _06804_ VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__o2bb2a_1
X_18966_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[8\] _11340_ _11387_
+ VGND VGND VPWR VPWR _11388_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17917_ _10038_ _10056_ _10420_ VGND VGND VPWR VPWR _10422_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_225_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18897_ _11308_ _11320_ VGND VGND VPWR VPWR _11321_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17848_ _10325_ _10326_ _10353_ VGND VGND VPWR VPWR _10355_ sky130_fd_sc_hd__nand3_1
XFILLER_0_191_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_233_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17779_ _10241_ _10243_ _10285_ VGND VGND VPWR VPWR _10287_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19518_ _11688_ _11700_ _01311_ _01310_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20790_ _02546_ _02542_ _02565_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19449_ _01281_ net236 _01245_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22460_ _04137_ _04141_ _04142_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__or3_1
XFILLER_0_29_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21411_ _03088_ _03096_ _03146_ VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22391_ _04030_ _04032_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24130_ clknet_leaf_118_clk _00663_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_21342_ _03077_ _03078_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24061_ clknet_leaf_45_clk _00594_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold620 top_inst.axis_out_inst.out_buff_data\[54\] VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__dlygate4sd3_1
X_21273_ top_inst.grid_inst.data_path_wires\[17\]\[3\] top_inst.grid_inst.data_path_wires\[17\]\[2\]
+ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__and4_1
Xhold631 _00204_ VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold642 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[13\] VGND
+ VGND VPWR VPWR net824 sky130_fd_sc_hd__dlygate4sd3_1
X_23012_ top_inst.axis_in_inst.inbuf_bus\[6\] _04588_ _04598_ _04590_ VGND VGND VPWR
+ VPWR _00980_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold653 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[2\] VGND
+ VGND VPWR VPWR net835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20224_ _01999_ _11163_ _02019_ _02006_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold664 top_inst.deskew_buff_inst.col_input\[8\] VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold675 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[12\] VGND
+ VGND VPWR VPWR net857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold686 top_inst.deskew_buff_inst.col_input\[94\] VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold697 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[25\] VGND
+ VGND VPWR VPWR net879 sky130_fd_sc_hd__dlygate4sd3_1
X_20155_ _01964_ _01965_ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20086_ _01890_ _01898_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__or2_1
XTAP_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_16
XTAP_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23914_ clknet_leaf_35_clk _00447_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[25\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23845_ clknet_leaf_96_clk _00378_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23776_ clknet_leaf_64_clk _00309_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11790_ net743 _04890_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__or2_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20988_ _02754_ _02755_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22727_ _04375_ _04368_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13460_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[7\] _05773_ VGND
+ VGND VPWR VPWR _06216_ sky130_fd_sc_hd__or2_1
X_22658_ _04329_ _04332_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12411_ net292 _05243_ _05249_ _05247_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21609_ _03272_ _03308_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13391_ _06136_ _06141_ _06163_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__a21o_1
X_22589_ _04262_ _04266_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__xor2_2
XFILLER_0_23_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_clk clknet_4_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_211_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15130_ _07779_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12342_ net650 _05204_ _05210_ _05208_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__o211a_1
X_24328_ clknet_leaf_5_clk _00861_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[18\]\[7\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_133_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15061_ top_inst.grid_inst.data_path_wires\[6\]\[1\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[6\]\[2\]
+ VGND VGND VPWR VPWR _07712_ sky130_fd_sc_hd__a22o_1
X_24259_ clknet_leaf_110_clk _00792_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_12273_ net879 _05169_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14012_ _06704_ _06729_ VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_1368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18820_ _11237_ _11245_ VGND VGND VPWR VPWR _11246_ sky130_fd_sc_hd__xor2_2
XFILLER_0_102_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18751_ _11135_ _11152_ _11132_ _11149_ VGND VGND VPWR VPWR _11180_ sky130_fd_sc_hd__nand4_1
XTAP_6185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15963_ _08532_ _08571_ VGND VGND VPWR VPWR _08573_ sky130_fd_sc_hd__and2_1
XFILLER_0_223_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_87_clk clknet_4_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_236_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17702_ top_inst.grid_inst.data_path_wires\[11\]\[0\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _10212_ sky130_fd_sc_hd__and2b_1
X_14914_ net1082 _07595_ VGND VGND VPWR VPWR _07596_ sky130_fd_sc_hd__and2_1
XTAP_5484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18682_ net706 _11116_ net167 VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__o21a_1
X_15894_ _08455_ _08454_ VGND VGND VPWR VPWR _08506_ sky130_fd_sc_hd__or2b_1
XTAP_5495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ _10111_ _10112_ _10144_ VGND VGND VPWR VPWR _10145_ sky130_fd_sc_hd__a21o_1
XFILLER_0_215_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14845_ _07087_ _07083_ _07090_ _07529_ VGND VGND VPWR VPWR _07530_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_192_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14776_ _07461_ _07462_ VGND VGND VPWR VPWR _07463_ sky130_fd_sc_hd__nand2_2
X_17564_ _10072_ _10078_ VGND VGND VPWR VPWR _10079_ sky130_fd_sc_hd__or2_1
X_11988_ _04994_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__clkbuf_4
X_19303_ _11701_ _11689_ VGND VGND VPWR VPWR _11702_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16515_ _09080_ _09048_ _09090_ VGND VGND VPWR VPWR _09092_ sky130_fd_sc_hd__nand3_1
X_13727_ _06427_ _06432_ _06471_ VGND VGND VPWR VPWR _06472_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_188_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17495_ _10025_ _07611_ _10026_ _10024_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19234_ _11514_ _11648_ VGND VGND VPWR VPWR _11649_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16446_ _09021_ _09024_ VGND VGND VPWR VPWR _09025_ sky130_fd_sc_hd__xor2_1
X_13658_ _06365_ _06360_ _06402_ _06404_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_144_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12609_ _05412_ _05421_ VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__xnor2_1
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16377_ _08870_ _08956_ _08957_ _08692_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__o211a_1
X_19165_ _11548_ _11544_ _11581_ _10957_ VGND VGND VPWR VPWR _11583_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13589_ _06193_ _06205_ _06334_ _06335_ VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__nand4_2
XFILLER_0_147_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk clknet_4_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15328_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[11\] _07845_ VGND
+ VGND VPWR VPWR _07973_ sky130_fd_sc_hd__xnor2_2
X_18116_ _10597_ _10057_ VGND VGND VPWR VPWR _10598_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19096_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[12\] _11340_ VGND
+ VGND VPWR VPWR _11515_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15259_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[9\] _07866_ VGND
+ VGND VPWR VPWR _07906_ sky130_fd_sc_hd__or2_1
X_18047_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[15\] _10367_ _10283_
+ VGND VGND VPWR VPWR _10548_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19998_ _01788_ _01815_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__xor2_1
XFILLER_0_226_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18949_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[7\] _11326_ _11371_
+ VGND VGND VPWR VPWR _11372_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_226_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_78_clk clknet_4_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_241_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21960_ _03279_ _03453_ _03673_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[27\]
+ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__a31o_1
XFILLER_0_193_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20911_ _05405_ _02681_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__nor2_1
X_21891_ _03311_ _03609_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23630_ clknet_leaf_102_clk net267 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_20842_ _02605_ _02606_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_230_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23561_ clknet_leaf_103_clk net701 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20773_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[17\] _02467_ VGND
+ VGND VPWR VPWR _02549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22512_ _04192_ _04169_ _04141_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23492_ clknet_leaf_140_clk net523 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[82\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22443_ _04092_ _04095_ _04097_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_49_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22374_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[11\] _03937_ _03938_
+ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24113_ clknet_leaf_16_clk _00646_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21325_ _02897_ _03062_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__xnor2_1
X_24044_ clknet_leaf_42_clk _00577_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold450 top_inst.axis_out_inst.out_buff_data\[11\] VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__dlygate4sd3_1
X_21256_ _02977_ _02973_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__or2b_1
XFILLER_0_241_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold461 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[1\] VGND VGND
+ VPWR VPWR net643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap180 _06934_ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__buf_1
Xhold472 top_inst.deskew_buff_inst.col_input\[111\] VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold483 top_inst.axis_out_inst.out_buff_data\[39\] VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__dlygate4sd3_1
X_20207_ _02007_ _11689_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__or2_1
Xhold494 top_inst.axis_out_inst.out_buff_data\[37\] VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21187_ _02868_ _02866_ _02885_ _02883_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__nand4_1
XFILLER_0_229_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20138_ net790 _01735_ _01949_ _01840_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__o211a_1
XTAP_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_69_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_16
XTAP_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20069_ _01882_ _01883_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__and2_1
X_12960_ _05268_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__clkbuf_8
XTAP_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ net868 _04951_ _04963_ _04955_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__o211a_1
XTAP_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12891_ _05335_ _05694_ _05695_ _05696_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__a31o_1
XFILLER_0_169_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1030 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[9\] _07281_ VGND
+ VGND VPWR VPWR _07320_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_174_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23828_ clknet_leaf_93_clk _00361_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11842_ net454 _04912_ _04924_ _04916_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__o211a_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _07234_ _07251_ _07252_ VGND VGND VPWR VPWR _07253_ sky130_fd_sc_hd__nand3_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _04859_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__clkbuf_4
X_23759_ clknet_leaf_122_clk net305 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _08833_ _08834_ _08881_ VGND VGND VPWR VPWR _08882_ sky130_fd_sc_hd__o21ba_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _06262_ VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__clkbuf_1
X_17280_ _09789_ _09788_ VGND VGND VPWR VPWR _09825_ sky130_fd_sc_hd__nand2_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14492_ net1125 _07152_ _07153_ VGND VGND VPWR VPWR _07186_ sky130_fd_sc_hd__nor3b_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16231_ _08806_ _08814_ VGND VGND VPWR VPWR _08815_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13443_ _05755_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16162_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[3\] _08728_ _08729_
+ VGND VGND VPWR VPWR _08748_ sky130_fd_sc_hd__a21bo_1
X_13374_ _05753_ _05770_ _05768_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15113_ _07755_ _07762_ VGND VGND VPWR VPWR _07763_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12325_ net943 _05191_ _05200_ _05195_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__o211a_1
X_16093_ _08688_ _08684_ VGND VGND VPWR VPWR _08689_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19921_ _01740_ _01741_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__nor2_2
X_15044_ _07610_ _07631_ VGND VGND VPWR VPWR _07696_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12256_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[18\] _05156_
+ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__or2_1
XFILLER_0_239_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19852_ net311 _01386_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__or2_1
XFILLER_0_236_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12187_ net799 _05115_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__or2_1
XFILLER_0_222_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18803_ _11205_ _11224_ VGND VGND VPWR VPWR _11229_ sky130_fd_sc_hd__nor2_1
X_19783_ _01486_ _01487_ _01607_ _01608_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__a211oi_2
X_16995_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[3\]
+ _09217_ VGND VGND VPWR VPWR _09549_ sky130_fd_sc_hd__and3_1
XFILLER_0_223_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18734_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[7\] _11150_ VGND
+ VGND VPWR VPWR _11166_ sky130_fd_sc_hd__or2_1
XTAP_5270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15946_ net1054 _05403_ VGND VGND VPWR VPWR _08556_ sky130_fd_sc_hd__nand2_1
XTAP_5281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_0_clk clknet_4_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_16
XTAP_5292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18665_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[16\] _10840_ _10791_
+ VGND VGND VPWR VPWR _11122_ sky130_fd_sc_hd__o21ba_1
XTAP_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15877_ _08487_ _08488_ VGND VGND VPWR VPWR _08489_ sky130_fd_sc_hd__xnor2_1
XTAP_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17616_ _10029_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[2\] VGND
+ VGND VPWR VPWR _10128_ sky130_fd_sc_hd__nand2_1
X_14828_ _07485_ _07475_ _07513_ VGND VGND VPWR VPWR _07514_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18596_ _11052_ _11055_ VGND VGND VPWR VPWR _11056_ sky130_fd_sc_hd__nor2_1
XFILLER_0_203_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17547_ net1041 _08183_ _10063_ _10049_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__o211a_1
X_14759_ _07404_ _07432_ _07431_ VGND VGND VPWR VPWR _07446_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_175_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17478_ _09661_ _10012_ VGND VGND VPWR VPWR _10013_ sky130_fd_sc_hd__and2_4
XFILLER_0_229_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19217_ _11621_ _11632_ VGND VGND VPWR VPWR _11633_ sky130_fd_sc_hd__xor2_1
XFILLER_0_116_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16429_ top_inst.grid_inst.data_path_wires\[8\]\[4\] top_inst.grid_inst.data_path_wires\[8\]\[5\]
+ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _09008_ sky130_fd_sc_hd__and4b_1
XFILLER_0_183_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19148_ _11479_ _11565_ VGND VGND VPWR VPWR _11566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19079_ _11495_ _11497_ VGND VGND VPWR VPWR _11499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21110_ top_inst.grid_inst.data_path_wires\[17\]\[3\] VGND VGND VPWR VPWR _02868_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22090_ _03707_ _03705_ _03684_ top_inst.grid_inst.data_path_wires\[18\]\[1\] VGND
+ VGND VPWR VPWR _03782_ sky130_fd_sc_hd__nand4_1
XFILLER_0_61_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21041_ _02760_ _02805_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__nor2_1
XFILLER_0_239_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22992_ top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[6\] _04583_ VGND
+ VGND VPWR VPWR _04587_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21943_ net561 _09804_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__or2_1
XFILLER_0_213_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_1252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21874_ _03568_ _03590_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__and2_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23613_ clknet_leaf_105_clk _00146_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20825_ _02596_ _02597_ _02473_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24593_ clknet_leaf_24_clk _01126_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_132_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23544_ clknet_leaf_130_clk _00077_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_20756_ _02514_ _02515_ _02531_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__or3_1
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23475_ clknet_leaf_136_clk _00008_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20687_ _02465_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__buf_2
XFILLER_0_68_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_443 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22426_ _04025_ _04074_ _04109_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_208_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22357_ _03999_ _04001_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12110_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[19\] _05076_
+ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21308_ _02871_ _02868_ _02891_ _02889_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__nand4_1
X_13090_ _05832_ _05870_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_237_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22288_ _03964_ _03966_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__nor2_1
X_24027_ clknet_leaf_48_clk _00560_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12041_ net782 _05031_ _05038_ _05035_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__o211a_1
Xhold280 top_inst.axis_out_inst.out_buff_data\[81\] VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__dlygate4sd3_1
X_21239_ _02972_ _02978_ VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_218_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold291 top_inst.axis_out_inst.out_buff_data\[101\] VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15800_ _08411_ _08413_ VGND VGND VPWR VPWR _08414_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_219_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16780_ _09337_ _09338_ VGND VGND VPWR VPWR _09339_ sky130_fd_sc_hd__nor2_1
X_13992_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[3\]
+ top_inst.grid_inst.data_path_wires\[3\]\[2\] top_inst.grid_inst.data_path_wires\[3\]\[1\]
+ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__nand4_1
XFILLER_0_189_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12943_ _05741_ _05735_ _05742_ _05743_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__o211a_1
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15731_ _08197_ _08346_ VGND VGND VPWR VPWR _08347_ sky130_fd_sc_hd__and2_1
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18450_ _10874_ _10913_ VGND VGND VPWR VPWR _10914_ sky130_fd_sc_hd__nand2_1
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ _05608_ _05679_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__nand2_1
XANTENNA_120 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _08163_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[2\] _08277_
+ _08278_ VGND VGND VPWR VPWR _08279_ sky130_fd_sc_hd__a22o_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _09913_ _09934_ _09939_ VGND VGND VPWR VPWR _09940_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14613_ _07302_ _07303_ VGND VGND VPWR VPWR _07304_ sky130_fd_sc_hd__xor2_1
X_11825_ net415 _04903_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__or2_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18381_ _10841_ _10845_ VGND VGND VPWR VPWR _10846_ sky130_fd_sc_hd__xor2_1
X_15593_ _08198_ _08192_ _08210_ VGND VGND VPWR VPWR _08213_ sky130_fd_sc_hd__and3_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _07070_ _07081_ VGND VGND VPWR VPWR _07236_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17332_ _09624_ _09873_ VGND VGND VPWR VPWR _09874_ sky130_fd_sc_hd__nor2_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11756_ net724 _04860_ _04872_ _04875_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__o211a_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14475_ _07162_ _07167_ _07168_ VGND VGND VPWR VPWR _07169_ sky130_fd_sc_hd__nand3_2
X_17263_ _09791_ _09797_ VGND VGND VPWR VPWR _09808_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19002_ _11382_ _11423_ VGND VGND VPWR VPWR _11424_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16214_ _08697_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[5\] _08664_
+ top_inst.grid_inst.data_path_wires\[8\]\[0\] VGND VGND VPWR VPWR _08798_ sky130_fd_sc_hd__nand4_2
X_13426_ _05177_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__clkbuf_4
X_17194_ _09741_ _09742_ VGND VGND VPWR VPWR _09743_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16145_ _08730_ _08731_ VGND VGND VPWR VPWR _08732_ sky130_fd_sc_hd__or2_2
XFILLER_0_52_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13357_ _06129_ _06114_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__and2b_1
XFILLER_0_52_986 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12308_ net909 _05178_ _05190_ _05182_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__o211a_1
X_16076_ top_inst.grid_inst.data_path_wires\[8\]\[6\] VGND VGND VPWR VPWR _08676_
+ sky130_fd_sc_hd__buf_2
X_13288_ _05751_ _06016_ _06017_ _05980_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19904_ _01721_ _01725_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__xor2_4
X_15027_ _07672_ _07679_ VGND VGND VPWR VPWR _07680_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12239_ _05044_ VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_209_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19835_ _01394_ _01524_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[16\]
+ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_224_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19766_ net596 _10616_ _01593_ _11714_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__o211a_1
X_16978_ _09454_ _09452_ _09491_ VGND VGND VPWR VPWR _09533_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 input_tdata[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_223_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18717_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _11154_ sky130_fd_sc_hd__buf_4
X_15929_ _08538_ _08539_ VGND VGND VPWR VPWR _08540_ sky130_fd_sc_hd__xnor2_2
X_19697_ _01524_ _01525_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_863 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18648_ _11099_ _11105_ VGND VGND VPWR VPWR _11106_ sky130_fd_sc_hd__xor2_1
XFILLER_0_231_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18579_ _11004_ _11003_ VGND VGND VPWR VPWR _11039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20610_ _02374_ _02376_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__or2b_1
XFILLER_0_117_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21590_ _03290_ _03293_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20541_ top_inst.grid_inst.data_path_wires\[16\]\[4\] _02020_ VGND VGND VPWR VPWR
+ _02324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23260_ net123 _04740_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20472_ _02224_ _02255_ _02256_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22211_ _03898_ _03899_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__nand2_1
X_23191_ net90 _04701_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22142_ _03820_ _03831_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22073_ _03707_ _03705_ top_inst.grid_inst.data_path_wires\[18\]\[1\] top_inst.grid_inst.data_path_wires\[18\]\[0\]
+ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__nand4_1
XTAP_6729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21024_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[25\] _02559_ _02789_
+ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22975_ top_inst.skew_buff_inst.row\[1\].output_reg\[6\] _04570_ VGND VGND VPWR VPWR
+ _04578_ sky130_fd_sc_hd__or2_1
XFILLER_0_214_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21926_ _03593_ _03642_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__and2_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21857_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[24\] _03421_ _03422_
+ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__a21oi_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20808_ _02581_ _02582_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__and2_1
X_24576_ clknet_leaf_142_clk _01109_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dfxtp_1
X_12590_ _05327_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__buf_8
XFILLER_0_136_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21788_ _03375_ _03496_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23527_ clknet_leaf_139_clk net649 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_955 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20739_ _02469_ _02499_ _02498_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14260_ _06926_ _06929_ _06927_ VGND VGND VPWR VPWR _06971_ sky130_fd_sc_hd__o21ba_1
X_23458_ net533 _04840_ _04851_ _04844_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13211_ _05945_ _05988_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22409_ _04092_ _04062_ _04064_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__o21bai_1
X_14191_ _06902_ _06889_ VGND VGND VPWR VPWR _06904_ sky130_fd_sc_hd__and2b_1
XFILLER_0_104_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23389_ net635 _04804_ _04814_ _04808_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13142_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[7\] _05326_ VGND
+ VGND VPWR VPWR _05922_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_237_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13073_ _05734_ _05770_ _05768_ _05738_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__a22o_1
X_17950_ _10413_ _10453_ VGND VGND VPWR VPWR _10454_ sky130_fd_sc_hd__nor2_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16901_ _09455_ _09456_ VGND VGND VPWR VPWR _09457_ sky130_fd_sc_hd__nand2_1
X_12024_ net315 _05018_ _05028_ _05022_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__o211a_1
X_17881_ _10377_ _10386_ VGND VGND VPWR VPWR _10387_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_228_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19620_ _01448_ _01449_ _01450_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__nand3_1
X_16832_ _09342_ _09344_ VGND VGND VPWR VPWR _09390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_228_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_232_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19551_ _01382_ _01383_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16763_ _08831_ _09322_ VGND VGND VPWR VPWR _09323_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13975_ _06618_ _06692_ _06693_ VGND VGND VPWR VPWR _06694_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_215_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18502_ _10963_ VGND VGND VPWR VPWR _10964_ sky130_fd_sc_hd__inv_2
XFILLER_0_232_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15714_ _08327_ _08328_ _08278_ _08280_ VGND VGND VPWR VPWR _08330_ sky130_fd_sc_hd__o211a_1
X_19482_ _01298_ net242 net190 _11703_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__a2bb2o_1
X_12926_ _05324_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__clkbuf_8
X_16694_ _09254_ _09255_ VGND VGND VPWR VPWR _09256_ sky130_fd_sc_hd__and2_1
XFILLER_0_186_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18433_ top_inst.grid_inst.data_path_wires\[12\]\[3\] _10614_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[6\]
+ top_inst.grid_inst.data_path_wires\[12\]\[4\] VGND VGND VPWR VPWR _10897_ sky130_fd_sc_hd__and4b_1
XFILLER_0_197_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15645_ _08260_ _08262_ VGND VGND VPWR VPWR _08263_ sky130_fd_sc_hd__xor2_1
X_12857_ _05636_ _05624_ _05663_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11808_ net576 _04898_ _04905_ _04902_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18364_ _10827_ _10829_ VGND VGND VPWR VPWR _10830_ sky130_fd_sc_hd__nand2_1
X_12788_ _05304_ _05567_ _05297_ _05302_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15576_ net1079 _08183_ _08196_ _08166_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__o211a_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _09853_ _09857_ VGND VGND VPWR VPWR _09858_ sky130_fd_sc_hd__xnor2_1
X_14527_ _07154_ _07185_ _07217_ _07218_ VGND VGND VPWR VPWR _07220_ sky130_fd_sc_hd__o22a_1
X_11739_ top_inst.axis_in_inst.inbuf_valid VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__inv_6
XFILLER_0_126_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18295_ top_inst.grid_inst.data_path_wires\[12\]\[3\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[3\] _10606_ VGND VGND
+ VPWR VPWR _10762_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17246_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[18\] _09628_ _09629_
+ VGND VGND VPWR VPWR _09792_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14458_ _07124_ _07126_ _07127_ _07123_ VGND VGND VPWR VPWR _07153_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13409_ net1035 _06169_ _06177_ _06179_ _06180_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__o221a_1
XFILLER_0_40_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14389_ top_inst.skew_buff_inst.row\[1\].output_reg\[7\] top_inst.axis_in_inst.inbuf_bus\[15\]
+ net212 VGND VGND VPWR VPWR _07089_ sky130_fd_sc_hd__mux2_2
X_17177_ _09678_ VGND VGND VPWR VPWR _09726_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16128_ _08714_ _08715_ VGND VGND VPWR VPWR _08716_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16059_ top_inst.grid_inst.data_path_wires\[8\]\[1\] VGND VGND VPWR VPWR _08664_
+ sky130_fd_sc_hd__buf_2
XFILLER_0_110_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19818_ _01642_ _01643_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__nor2_1
X_19749_ _01488_ _01575_ _01576_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__or3_1
XFILLER_0_155_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_237_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22760_ _04428_ _04429_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__nand2_2
XFILLER_0_91_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21711_ _03436_ _03437_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__and2_2
XFILLER_0_91_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22691_ _04284_ _04361_ _04363_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__a21o_1
XFILLER_0_220_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24430_ clknet_leaf_59_clk net882 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].output_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21642_ _03279_ _03353_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24361_ clknet_leaf_30_clk _00894_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[120\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_20 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21573_ _03302_ _03304_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__nor2_1
XFILLER_0_191_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_31 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_42 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23312_ net742 _04765_ _04771_ _04769_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__o211a_1
XANTENNA_53 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_209_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20524_ _02269_ _02307_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__xnor2_2
XANTENNA_64 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24292_ clknet_leaf_120_clk _00825_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_244_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_75 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_86 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23243_ net873 _04726_ _04732_ _04730_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__o211a_1
XANTENNA_97 _02707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20455_ _02238_ _02239_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__xor2_2
XFILLER_0_15_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23174_ net843 _04685_ _04693_ _04691_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20386_ top_inst.deskew_buff_inst.col_input\[38\] _11723_ _02171_ _02172_ VGND VGND
+ VPWR VPWR _02173_ sky130_fd_sc_hd__a22o_1
XFILLER_0_242_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22125_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[6\] _03814_ _03815_
+ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput160 net160 VGND VGND VPWR VPWR output_tdata[95] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22056_ _03742_ _03749_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__xnor2_1
XTAP_6559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21007_ _02749_ _02764_ _02773_ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__a21oi_2
XTAP_5858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_230_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13760_ _06499_ _06502_ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__and2_1
X_22958_ top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[7\] _04557_ VGND
+ VGND VPWR VPWR _04568_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12711_ _05476_ _05479_ _05520_ _05521_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__a211oi_2
X_21909_ _03595_ _03607_ _03625_ _01984_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13691_ _06335_ _06337_ _06386_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__and3_1
X_22889_ net728 _04522_ _04528_ _04524_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12642_ _05414_ _05453_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15430_ _08069_ _08070_ _07990_ _08071_ VGND VGND VPWR VPWR _08072_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_214_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24628_ clknet_leaf_24_clk _01161_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[104\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15361_ _07881_ _07954_ _07916_ VGND VGND VPWR VPWR _08005_ sky130_fd_sc_hd__o21ba_2
X_12573_ _05385_ _05386_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24559_ clknet_leaf_133_clk _01092_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_25_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17100_ _09650_ _09651_ VGND VGND VPWR VPWR _09652_ sky130_fd_sc_hd__nor2_2
XFILLER_0_0_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14312_ _07020_ _07021_ VGND VGND VPWR VPWR _07022_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15292_ _07935_ _07937_ VGND VGND VPWR VPWR _07938_ sky130_fd_sc_hd__xor2_1
X_18080_ net1002 _10563_ _10576_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_733 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17031_ _09573_ _09574_ VGND VGND VPWR VPWR _09584_ sky130_fd_sc_hd__nand2_1
X_14243_ _06869_ _06913_ _06954_ VGND VGND VPWR VPWR _06955_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14174_ _06848_ _06886_ _06887_ _06684_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13125_ _05750_ _05904_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__nand2_1
XFILLER_0_238_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18982_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[13\]\[3\]
+ _11135_ _11351_ VGND VGND VPWR VPWR _11404_ sky130_fd_sc_hd__o2bb2a_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _05822_ _05837_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__xnor2_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _10408_ _10437_ VGND VGND VPWR VPWR _10438_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_221_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12007_ net546 _05010_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17864_ _10040_ _10047_ _10336_ _10335_ _10038_ VGND VGND VPWR VPWR _10370_ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19603_ _01397_ _01400_ _01433_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__a21o_1
X_16815_ _09207_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[3\] _09201_
+ _09206_ VGND VGND VPWR VPWR _09373_ sky130_fd_sc_hd__and4_1
XFILLER_0_233_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17795_ _10298_ _10302_ VGND VGND VPWR VPWR _10303_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19534_ _01364_ _01365_ _01363_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__a21o_1
XFILLER_0_233_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1096 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16746_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[2\] _09202_ _09304_
+ _09305_ VGND VGND VPWR VPWR _09306_ sky130_fd_sc_hd__nand4_2
XFILLER_0_152_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13958_ _06676_ _06677_ VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__or2b_1
XFILLER_0_191_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12909_ _05655_ _05689_ _05687_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_198_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19465_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[6\] net231 _01263_
+ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__a21boi_1
X_16677_ _09232_ _09239_ VGND VGND VPWR VPWR _09240_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13889_ _06186_ _06192_ _06625_ _06446_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18416_ _10827_ _10829_ _10876_ VGND VGND VPWR VPWR _10880_ sky130_fd_sc_hd__a21o_1
XFILLER_0_232_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15628_ _08239_ _08244_ VGND VGND VPWR VPWR _08246_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19396_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[5\] _01230_ _01231_
+ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18347_ _10810_ _10812_ VGND VGND VPWR VPWR _10813_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15559_ _05335_ VGND VGND VPWR VPWR _08181_ sky130_fd_sc_hd__buf_6
XFILLER_0_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18278_ _10656_ _10678_ _10703_ _10707_ VGND VGND VPWR VPWR _10746_ sky130_fd_sc_hd__o31a_1
XFILLER_0_142_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17229_ _09774_ _09775_ VGND VGND VPWR VPWR _09776_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold802 _00975_ VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold813 top_inst.axis_in_inst.inbuf_bus\[13\] VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__dlygate4sd3_1
X_20240_ _02030_ _02031_ _02024_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__a21oi_1
Xhold824 top_inst.axis_in_inst.inbuf_bus\[31\] VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold835 top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[0\] VGND VGND
+ VPWR VPWR net1017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold846 top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[27\] VGND VGND
+ VPWR VPWR net1028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_243_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold857 top_inst.axis_in_inst.inbuf_bus\[26\] VGND VGND VPWR VPWR net1039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold868 top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[21\] VGND VGND
+ VPWR VPWR net1050 sky130_fd_sc_hd__dlygate4sd3_1
X_20171_ _01975_ _01980_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold879 top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[9\] VGND VGND
+ VPWR VPWR net1061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23930_ clknet_leaf_75_clk _00463_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23861_ clknet_leaf_77_clk _00394_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_93_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22812_ _07707_ _04478_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23792_ clknet_leaf_71_clk _00325_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22743_ _04412_ _04413_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22674_ _04346_ _04347_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__and2b_1
XFILLER_0_133_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24413_ clknet_leaf_56_clk net591 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21625_ _03352_ _03354_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_164_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24344_ clknet_leaf_8_clk _00877_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[103\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21556_ top_inst.grid_inst.data_path_wires\[17\]\[6\] _02897_ VGND VGND VPWR VPWR
+ _03288_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_106_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_244_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20507_ _02241_ _02288_ _02289_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__nor3_1
XFILLER_0_244_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24275_ clknet_leaf_11_clk _00808_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[17\]\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_21487_ _03171_ _03179_ _03220_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_132_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23226_ net731 _04713_ _04722_ _04717_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20438_ _02177_ _02183_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__and2b_1
XFILLER_0_244_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23157_ net75 _04672_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__or2_1
XTAP_6301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20369_ _02152_ _02153_ _02154_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__a21o_1
XTAP_6312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22108_ _03751_ _03773_ _03799_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__o21ai_1
XTAP_6334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23088_ net1113 _04602_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__or2_1
XTAP_5600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14930_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[27\] _07576_ VGND
+ VGND VPWR VPWR _07604_ sky130_fd_sc_hd__and2_1
XTAP_5633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22039_ _03732_ _03733_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__and2_1
XTAP_6389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14861_ _07544_ _07545_ VGND VGND VPWR VPWR _07546_ sky130_fd_sc_hd__nand2_1
XFILLER_0_215_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600_ _09156_ _09173_ VGND VGND VPWR VPWR _09174_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ _06554_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17580_ _10091_ _10092_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[3\]
+ VGND VGND VPWR VPWR _10094_ sky130_fd_sc_hd__a21oi_1
X_14792_ _07445_ _07478_ VGND VGND VPWR VPWR _07479_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_203_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16531_ _09105_ _09107_ VGND VGND VPWR VPWR _09108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13743_ _06193_ _06214_ _06485_ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19250_ _11645_ _11651_ _11653_ VGND VGND VPWR VPWR _11664_ sky130_fd_sc_hd__o21a_1
X_16462_ _08679_ _08695_ VGND VGND VPWR VPWR _09040_ sky130_fd_sc_hd__nand2_2
XFILLER_0_35_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13674_ _06418_ _06419_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_1302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18201_ _10581_ _10602_ VGND VGND VPWR VPWR _10671_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15413_ _08013_ _08015_ VGND VGND VPWR VPWR _08056_ sky130_fd_sc_hd__or2b_1
XPHY_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12625_ _05435_ _05436_ _05407_ _05398_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__o211a_1
XFILLER_0_182_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19181_ _11147_ _11161_ VGND VGND VPWR VPWR _11598_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16393_ _08971_ _08959_ VGND VGND VPWR VPWR _08973_ sky130_fd_sc_hd__and2b_1
XPHY_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18132_ _10606_ _10607_ _10609_ _10594_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__o211a_1
X_12556_ _05356_ _05370_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15344_ _05632_ _07988_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18063_ _05313_ VGND VGND VPWR VPWR _10563_ sky130_fd_sc_hd__clkbuf_4
X_12487_ _05269_ _05306_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15275_ _07908_ _07920_ VGND VGND VPWR VPWR _07921_ sky130_fd_sc_hd__and2b_1
XFILLER_0_123_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17014_ _09565_ _09566_ _09548_ VGND VGND VPWR VPWR _09568_ sky130_fd_sc_hd__a21oi_1
Xhold109 _01160_ VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__dlygate4sd3_1
X_14226_ _06895_ _06896_ VGND VGND VPWR VPWR _06938_ sky130_fd_sc_hd__or2b_1
XFILLER_0_238_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14157_ _06869_ _06870_ VGND VGND VPWR VPWR _06871_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13108_ _05856_ _05861_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__nor2_1
X_14088_ _06801_ _06802_ _05633_ VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__a21o_1
X_18965_ _11339_ VGND VGND VPWR VPWR _11387_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13039_ _05821_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__clkbuf_1
X_17916_ _10037_ _10056_ _10420_ VGND VGND VPWR VPWR _10421_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18896_ _11313_ _11319_ VGND VGND VPWR VPWR _11320_ sky130_fd_sc_hd__xor2_1
XFILLER_0_206_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17847_ _10325_ _10326_ _10353_ VGND VGND VPWR VPWR _10354_ sky130_fd_sc_hd__a21o_1
XFILLER_0_240_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17778_ _10241_ _10243_ _10285_ VGND VGND VPWR VPWR _10286_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19517_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[7\] _01302_ _01301_
+ _11684_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__a22o_1
X_16729_ _09259_ _09262_ VGND VGND VPWR VPWR _09290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19448_ _01245_ _01281_ _01282_ VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_232_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19379_ _01213_ _01214_ _01212_ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21410_ _03093_ _03095_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__and2_1
XFILLER_0_228_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22390_ _04025_ _04074_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21341_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[1\] _02882_ top_inst.grid_inst.data_path_wires\[17\]\[7\]
+ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_170_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24060_ clknet_leaf_45_clk _00593_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold610 _00096_ VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__dlygate4sd3_1
X_21272_ top_inst.grid_inst.data_path_wires\[17\]\[2\] _02891_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[3\]
+ top_inst.grid_inst.data_path_wires\[17\]\[3\] VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_13_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold621 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[8\] VGND
+ VGND VPWR VPWR net803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23011_ net1063 _04596_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold632 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[24\] VGND
+ VGND VPWR VPWR net814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold643 top_inst.deskew_buff_inst.col_input\[22\] VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__dlygate4sd3_1
X_20223_ _02018_ _11689_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold654 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[21\] VGND
+ VGND VPWR VPWR net836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold665 _00207_ VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[2\] VGND
+ VGND VPWR VPWR net858 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold687 top_inst.deskew_buff_inst.col_input\[60\] VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__dlygate4sd3_1
X_20154_ _01944_ _01945_ _01963_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__o21bai_1
Xhold698 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[7\] VGND
+ VGND VPWR VPWR net880 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20085_ _01890_ _01898_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__nand2_1
XTAP_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23913_ clknet_leaf_33_clk _00446_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23844_ clknet_leaf_96_clk _00377_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23775_ clknet_leaf_63_clk _00308_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20987_ _02725_ _02740_ _02753_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__nand3_1
XFILLER_0_71_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22726_ _04386_ _04397_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22657_ _04331_ _04327_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__xor2_2
XFILLER_0_211_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12410_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[20\] _05248_
+ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__or2_1
XFILLER_0_193_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21608_ _03305_ _03338_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__xor2_1
XFILLER_0_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13390_ _06161_ _06162_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22588_ _04264_ _04265_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__and2b_1
XFILLER_0_129_1016 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12341_ net333 _05209_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21539_ _03239_ _03271_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__xor2_2
X_24327_ clknet_leaf_5_clk _00860_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[18\]\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_209_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15060_ _07606_ _07637_ VGND VGND VPWR VPWR _07711_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24258_ clknet_leaf_110_clk _00791_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_12272_ net786 _05164_ _05170_ _05168_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14011_ _06727_ _06728_ VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23209_ net665 _04700_ _04712_ _04704_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24189_ clknet_leaf_47_clk _00722_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_219_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18750_ _11152_ _11132_ _11149_ _11135_ VGND VGND VPWR VPWR _11179_ sky130_fd_sc_hd__a22o_1
XTAP_6175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15962_ _08532_ _08571_ VGND VGND VPWR VPWR _08572_ sky130_fd_sc_hd__nor2_1
XTAP_5441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17701_ top_inst.grid_inst.data_path_wires\[11\]\[1\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _10211_ sky130_fd_sc_hd__nand2_1
XTAP_5463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14913_ _05633_ VGND VGND VPWR VPWR _07595_ sky130_fd_sc_hd__buf_8
XFILLER_0_222_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18681_ net1028 _11116_ net167 VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__o21a_1
XFILLER_0_236_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15893_ _08503_ _08504_ VGND VGND VPWR VPWR _08505_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_215_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17632_ _10089_ _10110_ VGND VGND VPWR VPWR _10144_ sky130_fd_sc_hd__nor2_1
X_14844_ _07459_ _07499_ _07497_ VGND VGND VPWR VPWR _07529_ sky130_fd_sc_hd__o21a_1
XTAP_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_926 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17563_ _10076_ _10077_ VGND VGND VPWR VPWR _10078_ sky130_fd_sc_hd__xor2_1
X_14775_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[7\] _07416_ _07085_
+ _07087_ VGND VGND VPWR VPWR _07462_ sky130_fd_sc_hd__a22o_1
X_11987_ net1108 _04996_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19302_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _11701_ sky130_fd_sc_hd__buf_2
XFILLER_0_187_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16514_ _09080_ _09048_ _09090_ VGND VGND VPWR VPWR _09091_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13726_ _06426_ _06423_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__and2b_1
X_17494_ _05736_ _09192_ VGND VGND VPWR VPWR _10026_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19233_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[16\] _11469_ VGND
+ VGND VPWR VPWR _11648_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16445_ _09022_ _09023_ VGND VGND VPWR VPWR _09024_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13657_ _05325_ VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_184_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12608_ _05415_ _05420_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__xor2_1
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19164_ _11548_ _11544_ _11581_ VGND VGND VPWR VPWR _11582_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16376_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[9\] _07866_ VGND
+ VGND VPWR VPWR _08957_ sky130_fd_sc_hd__or2_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13588_ top_inst.grid_inst.data_path_wires\[2\]\[5\] _06205_ _06334_ _06335_ VGND
+ VGND VPWR VPWR _06336_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18115_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _10597_ sky130_fd_sc_hd__clkbuf_4
X_15327_ _07624_ _07631_ _07917_ _07916_ _07622_ VGND VGND VPWR VPWR _07972_ sky130_fd_sc_hd__a32o_1
XFILLER_0_26_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19095_ _11513_ VGND VGND VPWR VPWR _11514_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12539_ _05353_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__buf_8
XFILLER_0_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18046_ _10545_ _10498_ VGND VGND VPWR VPWR _10547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15258_ _07868_ _07904_ VGND VGND VPWR VPWR _07905_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14209_ _06919_ _06920_ _06404_ VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__a21o_1
XFILLER_0_160_1338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15189_ _07831_ _07836_ VGND VGND VPWR VPWR _07837_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_239_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19997_ _01813_ _01814_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__nor2_1
XFILLER_0_238_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18948_ _11325_ _11324_ VGND VGND VPWR VPWR _11371_ sky130_fd_sc_hd__and2b_1
XFILLER_0_236_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18879_ top_inst.grid_inst.data_path_wires\[13\]\[7\] top_inst.grid_inst.data_path_wires\[13\]\[6\]
+ _11152_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _11303_ sky130_fd_sc_hd__nand4_1
XFILLER_0_241_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_234_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20910_ _02656_ _02680_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21890_ _05312_ _03595_ _03606_ _03607_ _03608_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__a41o_1
XFILLER_0_179_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20841_ _02581_ _02608_ _02607_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23560_ clknet_leaf_100_clk _00093_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20772_ _02518_ _02525_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22511_ _04025_ _04136_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__or2_2
XFILLER_0_130_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23491_ clknet_leaf_139_clk _00024_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[81\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22442_ _04114_ _04093_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__or2b_1
XFILLER_0_29_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22373_ _04016_ _04019_ _04057_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_206_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24112_ clknet_leaf_16_clk _00645_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21324_ _03060_ _03061_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24043_ clknet_leaf_42_clk _00576_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[19\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold440 top_inst.axis_out_inst.out_buff_data\[65\] VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__dlygate4sd3_1
X_21255_ _02981_ _02983_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold451 top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[7\] VGND VGND
+ VPWR VPWR net633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 _00951_ VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap170 _09313_ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
Xhold473 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[2\] VGND VGND
+ VPWR VPWR net655 sky130_fd_sc_hd__dlygate4sd3_1
X_20206_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _02007_ sky130_fd_sc_hd__clkbuf_4
Xmax_cap181 _06494_ VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__buf_1
Xhold484 top_inst.deskew_buff_inst.col_input\[125\] VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold495 top_inst.axis_out_inst.out_buff_data\[2\] VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__dlygate4sd3_1
X_21186_ _02866_ _02885_ _02882_ _02868_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__a22o_1
XFILLER_0_217_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20137_ _01932_ _01947_ _01948_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20068_ _01857_ _01881_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__or2_1
XTAP_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ net689 _04956_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__or2_1
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[13\] _05326_ VGND
+ VGND VPWR VPWR _05696_ sky130_fd_sc_hd__and2_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_1042 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23827_ clknet_leaf_93_clk _00360_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_11841_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[0\] _04917_
+ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__or2_1
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14560_ _07249_ _07250_ _07235_ VGND VGND VPWR VPWR _07252_ sky130_fd_sc_hd__a21o_1
XFILLER_0_166_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11772_ net888 _04860_ _04884_ _04875_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__o211a_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23758_ clknet_leaf_121_clk _00291_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13511_ _05886_ _06261_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__and2_1
X_22709_ _04380_ _04381_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_1096 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14491_ _07183_ _07184_ VGND VGND VPWR VPWR _07185_ sky130_fd_sc_hd__or2_2
XFILLER_0_166_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23689_ clknet_leaf_119_clk _00222_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16230_ _08807_ _08813_ VGND VGND VPWR VPWR _08814_ sky130_fd_sc_hd__xnor2_1
X_13442_ _06184_ _05756_ _06203_ _06183_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16161_ _08725_ _08746_ VGND VGND VPWR VPWR _08747_ sky130_fd_sc_hd__xnor2_2
X_13373_ _06099_ _06128_ _06145_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15112_ _07760_ _07761_ VGND VGND VPWR VPWR _07762_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12324_ net505 _05196_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__or2_1
X_16092_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _08688_ sky130_fd_sc_hd__buf_4
XFILLER_0_133_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19920_ _01561_ _01739_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15043_ _07693_ _07694_ VGND VGND VPWR VPWR _07695_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12255_ net968 _05151_ _05160_ _05155_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19851_ _01674_ _01675_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__and2_1
X_12186_ net759 _05110_ _05120_ _05114_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__o211a_1
X_18802_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[4\] _10364_ _11226_
+ _11227_ _11228_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__o221a_1
X_19782_ _01607_ _01608_ _01486_ _01487_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16994_ _09544_ _09547_ VGND VGND VPWR VPWR _09548_ sky130_fd_sc_hd__xor2_1
XFILLER_0_236_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18733_ _11145_ _11163_ _11165_ _11160_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__o211a_1
XTAP_5260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15945_ _08555_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18664_ _11100_ _11104_ VGND VGND VPWR VPWR _11121_ sky130_fd_sc_hd__nand2_1
XFILLER_0_222_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15876_ _08149_ _08167_ VGND VGND VPWR VPWR _08488_ sky130_fd_sc_hd__nand2_1
XTAP_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17615_ _10022_ _10054_ VGND VGND VPWR VPWR _10127_ sky130_fd_sc_hd__nand2_1
X_14827_ _07511_ _07512_ VGND VGND VPWR VPWR _07513_ sky130_fd_sc_hd__nor2_1
XFILLER_0_231_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18595_ _10612_ _11053_ _11014_ _11054_ VGND VGND VPWR VPWR _11055_ sky130_fd_sc_hd__a22oi_2
XTAP_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17546_ _10061_ _10062_ _08181_ VGND VGND VPWR VPWR _10063_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14758_ _07434_ _07435_ VGND VGND VPWR VPWR _07445_ sky130_fd_sc_hd__or2b_1
XFILLER_0_188_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13709_ top_inst.grid_inst.data_path_wires\[2\]\[5\] _06212_ VGND VGND VPWR VPWR
+ _06454_ sky130_fd_sc_hd__nand2_1
X_17477_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[30\] _10010_ _08307_
+ VGND VGND VPWR VPWR _10012_ sky130_fd_sc_hd__mux2_2
X_14689_ _07078_ VGND VGND VPWR VPWR _07378_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19216_ _11630_ _11631_ VGND VGND VPWR VPWR _11632_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16428_ _08932_ _09006_ VGND VGND VPWR VPWR _09007_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19147_ _11563_ _11564_ VGND VGND VPWR VPWR _11565_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16359_ _08885_ _08887_ _08939_ VGND VGND VPWR VPWR _08940_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19078_ _11495_ _11497_ VGND VGND VPWR VPWR _11498_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_1211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18029_ _10523_ _10530_ VGND VGND VPWR VPWR _10531_ sky130_fd_sc_hd__xor2_1
XFILLER_0_199_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21040_ _02779_ _02801_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__or2b_1
XFILLER_0_22_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22991_ net995 _04575_ _04586_ _04577_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__o211a_1
XFILLER_0_242_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21942_ _03648_ _03657_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21873_ net953 _03528_ _03591_ _03592_ _02962_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__o221a_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23612_ clknet_leaf_105_clk _00145_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_20824_ _02466_ _02596_ _02597_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24592_ clknet_leaf_22_clk _01125_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_38_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23543_ clknet_leaf_130_clk _00076_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_20755_ _02514_ _02515_ _02531_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_92_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23474_ clknet_leaf_134_clk net626 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20686_ _02004_ _02018_ _02438_ _02227_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__a31o_2
XFILLER_0_92_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22425_ _04071_ _04073_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__and2_1
XFILLER_0_162_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22356_ _04015_ _04041_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__xor2_2
XFILLER_0_131_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21307_ top_inst.grid_inst.data_path_wires\[17\]\[3\] _02891_ _02889_ top_inst.grid_inst.data_path_wires\[17\]\[4\]
+ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22287_ net964 _03528_ _03973_ _03974_ _02962_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__o221a_1
XFILLER_0_206_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24026_ clknet_leaf_48_clk _00559_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12040_ net469 _05036_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_1328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold270 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[5\] VGND
+ VGND VPWR VPWR net452 sky130_fd_sc_hd__dlygate4sd3_1
X_21238_ _02973_ _02977_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_236_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold281 top_inst.axis_out_inst.out_buff_data\[3\] VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold292 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[22\] VGND
+ VGND VPWR VPWR net474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21169_ _02866_ _02864_ _02885_ _02883_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__nand4_1
XFILLER_0_244_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_219_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13991_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[3\]\[2\]
+ top_inst.grid_inst.data_path_wires\[3\]\[1\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[4\]
+ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15730_ _08344_ _08345_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[7\]
+ _07816_ VGND VGND VPWR VPWR _08346_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_204_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12942_ _05260_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ top_inst.grid_inst.data_path_wires\[7\]\[3\] _08139_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _08278_ sky130_fd_sc_hd__nand4_2
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12873_ _05677_ _05678_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__and2_1
XANTENNA_110 _05313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_121 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17400_ _09937_ _09938_ VGND VGND VPWR VPWR _09939_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _07251_ _07253_ VGND VGND VPWR VPWR _07303_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ net889 _04912_ _04914_ _04902_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__o211a_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ _10843_ _10844_ VGND VGND VPWR VPWR _10845_ sky130_fd_sc_hd__nor2_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _08211_ VGND VGND VPWR VPWR _08212_ sky130_fd_sc_hd__inv_2
XFILLER_0_200_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[23\] _09631_ VGND
+ VGND VPWR VPWR _09873_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _07202_ _07203_ _07206_ VGND VGND VPWR VPWR _07235_ sky130_fd_sc_hd__and3_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _04874_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__buf_4
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17262_ _09798_ _09799_ VGND VGND VPWR VPWR _09807_ sky130_fd_sc_hd__and2b_1
XFILLER_0_153_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14474_ _07165_ _07166_ _07146_ _07148_ VGND VGND VPWR VPWR _07168_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_125_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19001_ _11383_ _11422_ VGND VGND VPWR VPWR _11423_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16213_ _08695_ _08664_ top_inst.grid_inst.data_path_wires\[8\]\[0\] _08697_ VGND
+ VGND VPWR VPWR _08797_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13425_ _05746_ _05256_ _06191_ _06183_ VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17193_ _09712_ _09740_ VGND VGND VPWR VPWR _09742_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16144_ _08728_ _08729_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[3\]
+ VGND VGND VPWR VPWR _08731_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13356_ _06114_ _06129_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12307_ net568 _05183_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__or2_1
X_16075_ _08147_ _08663_ _08675_ _08666_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__o211a_1
X_13287_ _06061_ _06062_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_886 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19903_ _01723_ _01724_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__and2b_1
X_15026_ _07677_ _07678_ VGND VGND VPWR VPWR _07679_ sky130_fd_sc_hd__xnor2_1
X_12238_ net426 _05137_ _05150_ _05141_ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_209_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19834_ _01352_ _01353_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[16\]
+ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__or3b_1
X_12169_ net317 _05102_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__or2_1
XFILLER_0_208_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16977_ _09497_ _09531_ VGND VGND VPWR VPWR _09532_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19765_ _05317_ _01592_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 input_tdata[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
XFILLER_0_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18716_ _11132_ _10607_ _11153_ _11137_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15928_ _08496_ _08502_ _08495_ VGND VGND VPWR VPWR _08539_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19696_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[11\] _01480_ VGND
+ VGND VPWR VPWR _01525_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18647_ _11100_ _11104_ VGND VGND VPWR VPWR _11105_ sky130_fd_sc_hd__xor2_1
XFILLER_0_210_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15859_ _08469_ _08471_ VGND VGND VPWR VPWR _08472_ sky130_fd_sc_hd__nand2_1
XFILLER_0_232_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18578_ net1085 _10364_ _11037_ _11038_ _09886_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__o221a_1
XFILLER_0_188_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17529_ _10050_ _09199_ VGND VGND VPWR VPWR _10051_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20540_ _02315_ _02322_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__xor2_1
XFILLER_0_28_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20471_ _02253_ _02254_ _02202_ _02225_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__a211o_1
XFILLER_0_229_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22210_ _03690_ _03707_ _03688_ _03705_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__nand4_1
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23190_ net492 _04700_ _04702_ _04691_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22141_ _03820_ _03831_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22072_ _03703_ _03684_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__nand2_2
XTAP_6719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21023_ _02473_ _02788_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1084 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22974_ net881 _04575_ _04576_ _04577_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21925_ _03606_ _03607_ _03625_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__and3_1
XFILLER_0_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24644_ clknet_leaf_21_clk net442 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[120\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21856_ _03574_ _03575_ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__nand2_2
XFILLER_0_78_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20807_ _02517_ _02573_ _02580_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__nand3_1
XFILLER_0_93_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24575_ clknet_leaf_142_clk _01108_ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dfxtp_2
X_21787_ _03469_ _03486_ _03506_ _03509_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_136_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23526_ clknet_leaf_1_clk net887 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20738_ _02495_ _02505_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23457_ top_inst.axis_out_inst.out_buff_data\[116\] _04864_ VGND VGND VPWR VPWR _04851_
+ sky130_fd_sc_hd__or2_1
X_20669_ _02411_ _02413_ _02448_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_243_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13210_ _05987_ _05938_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__nor2_1
X_22408_ _04061_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14190_ _06889_ _06902_ VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__and2b_1
XFILLER_0_150_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23388_ net57 _04805_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13141_ net169 _05881_ _05919_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22339_ _03950_ _04024_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_108_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13072_ _05823_ _05828_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_1163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16900_ _09414_ _09421_ VGND VGND VPWR VPWR _09456_ sky130_fd_sc_hd__or2b_1
X_12023_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[14\] _05023_
+ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__or2_1
X_24009_ clknet_leaf_47_clk _00542_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_17880_ _10384_ _10385_ VGND VGND VPWR VPWR _10386_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16831_ _09386_ _09387_ _09369_ VGND VGND VPWR VPWR _09389_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19550_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[7\] _01334_ _01333_
+ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__a21o_1
X_16762_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[5\] _09321_ _08307_
+ VGND VGND VPWR VPWR _09322_ sky130_fd_sc_hd__mux2_1
X_13974_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[3\]\[1\]
+ top_inst.grid_inst.data_path_wires\[3\]\[0\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[4\]
+ VGND VGND VPWR VPWR _06693_ sky130_fd_sc_hd__a22o_1
XFILLER_0_232_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18501_ _10924_ _10929_ _10927_ VGND VGND VPWR VPWR _10963_ sky130_fd_sc_hd__a21o_1
XFILLER_0_219_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15713_ _08278_ _08280_ _08327_ _08328_ VGND VGND VPWR VPWR _08329_ sky130_fd_sc_hd__a211oi_1
X_12925_ _05724_ _05728_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__xnor2_1
X_19481_ _01297_ _01314_ _11676_ net189 VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__or4b_4
X_16693_ _09203_ _09198_ _09186_ _09192_ VGND VGND VPWR VPWR _09255_ sky130_fd_sc_hd__nand4_2
XFILLER_0_232_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18432_ _10589_ _10610_ VGND VGND VPWR VPWR _10896_ sky130_fd_sc_hd__nand2_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15644_ _08211_ _08233_ _08261_ VGND VGND VPWR VPWR _08262_ sky130_fd_sc_hd__o21a_1
X_12856_ _05616_ _05662_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11807_ net462 _04903_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__or2_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _10781_ _10782_ _10828_ VGND VGND VPWR VPWR _10829_ sky130_fd_sc_hd__a21o_1
XFILLER_0_201_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15575_ _08194_ _08195_ _06682_ VGND VGND VPWR VPWR _08196_ sky130_fd_sc_hd__a21o_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _05561_ _05595_ _05440_ VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _09855_ _09856_ VGND VGND VPWR VPWR _09857_ sky130_fd_sc_hd__xor2_1
XFILLER_0_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14526_ _07154_ _07185_ _07217_ _07218_ VGND VGND VPWR VPWR _07219_ sky130_fd_sc_hd__nor4_4
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18294_ _10727_ _10732_ VGND VGND VPWR VPWR _10761_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11738_ _04859_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__buf_4
XFILLER_0_113_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17245_ _09625_ _09772_ _09790_ VGND VGND VPWR VPWR _09791_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14457_ _07143_ _07144_ _07150_ VGND VGND VPWR VPWR _07152_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13408_ _04874_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__clkbuf_16
X_17176_ _09703_ _09705_ _09724_ VGND VGND VPWR VPWR _09725_ sky130_fd_sc_hd__a21o_1
X_14388_ _05290_ _07086_ _07088_ _06684_ VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16127_ _08704_ _08705_ VGND VGND VPWR VPWR _08715_ sky130_fd_sc_hd__nand2_1
X_13339_ _06097_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16058_ _05177_ VGND VGND VPWR VPWR _08663_ sky130_fd_sc_hd__buf_4
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15009_ _07655_ _07661_ VGND VGND VPWR VPWR _07663_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19817_ _01629_ _01617_ _01641_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__and3_1
XFILLER_0_224_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19748_ _01573_ _01574_ _01570_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_1180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19679_ _01434_ _01461_ _01460_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21710_ _03414_ _03435_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__or2_1
X_22690_ _04325_ _04360_ _04357_ _04362_ _04356_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__a32o_1
XFILLER_0_154_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21641_ _03362_ _03364_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24360_ clknet_leaf_30_clk _00893_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[119\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21572_ _03243_ _03267_ _03303_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_10 top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[0\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_21 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_32 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_43 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23311_ net147 _04766_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__or2_1
X_20523_ _02305_ _02306_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__xnor2_2
XANTENNA_54 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24291_ clknet_leaf_120_clk _00824_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_65 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_209_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_76 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_87 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23242_ net114 _04727_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__or2_1
XANTENNA_98 _02707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20454_ _01995_ _02018_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23173_ net81 _04687_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__or2_1
X_20385_ _02136_ _02170_ _05399_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22124_ top_inst.grid_inst.data_path_wires\[18\]\[6\] top_inst.grid_inst.data_path_wires\[18\]\[5\]
+ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[1\] _03697_ VGND VGND
+ VPWR VPWR _03815_ sky130_fd_sc_hd__nand4_1
XFILLER_0_63_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput150 net150 VGND VGND VPWR VPWR output_tdata[86] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_219_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput161 net161 VGND VGND VPWR VPWR output_tdata[96] sky130_fd_sc_hd__clkbuf_4
XTAP_6516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22055_ _03747_ _03748_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__xnor2_2
XTAP_6549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21006_ _02771_ _02772_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__xnor2_1
XTAP_5837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_242_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22957_ net621 _04562_ _04567_ _04564_ VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_214_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12710_ _05518_ _05519_ _05472_ _05474_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__o211a_1
X_21908_ _03595_ _03607_ _03625_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13690_ _06433_ _06435_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__xnor2_1
X_22888_ net578 _04517_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__or2_1
XFILLER_0_179_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_1416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12641_ _05451_ _05452_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__xor2_1
XFILLER_0_194_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24627_ clknet_leaf_23_clk net291 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[103\]
+ sky130_fd_sc_hd__dfxtp_1
X_21839_ _03555_ _03559_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15360_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[11\] _07924_ _07844_
+ VGND VGND VPWR VPWR _08004_ sky130_fd_sc_hd__a21o_1
X_12572_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[1\] _05292_ _05296_
+ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _05386_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_136_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24558_ clknet_leaf_135_clk _01091_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_38_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14311_ _06989_ _06992_ _06987_ VGND VGND VPWR VPWR _07021_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23509_ clknet_leaf_136_clk net314 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15291_ _07896_ _07897_ _07936_ VGND VGND VPWR VPWR _07937_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24489_ clknet_leaf_45_clk net332 VGND VGND VPWR VPWR top_inst.valid_pipe\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17030_ _09533_ _09579_ _09580_ _09409_ _09582_ VGND VGND VPWR VPWR _09583_ sky130_fd_sc_hd__o221a_4
XFILLER_0_150_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14242_ _06910_ _06912_ VGND VGND VPWR VPWR _06954_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_499 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14173_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[9\] _06168_ VGND
+ VGND VPWR VPWR _06887_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13124_ top_inst.grid_inst.data_path_wires\[1\]\[7\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _05904_ sky130_fd_sc_hd__and3_1
X_18981_ top_inst.grid_inst.data_path_wires\[13\]\[2\] top_inst.grid_inst.data_path_wires\[13\]\[3\]
+ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _11403_ sky130_fd_sc_hd__and4b_1
XFILLER_0_238_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13055_ _05829_ _05836_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__xor2_2
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17932_ _10435_ _10436_ VGND VGND VPWR VPWR _10437_ sky130_fd_sc_hd__nand2_1
X_12006_ _04911_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__buf_2
XFILLER_0_139_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17863_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[11\] _10236_ VGND
+ VGND VPWR VPWR _10369_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_205_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19602_ _01399_ _01398_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16814_ _09207_ _09202_ _09206_ _09203_ VGND VGND VPWR VPWR _09372_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_89_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17794_ _10299_ _10301_ VGND VGND VPWR VPWR _10302_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1039 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16745_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[3\]
+ net1119 net225 VGND VGND VPWR VPWR _09305_ sky130_fd_sc_hd__nand4_4
X_19533_ _01363_ _01364_ _01365_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__nand3_1
XFILLER_0_117_1316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13957_ _06673_ _06674_ _06675_ _06671_ VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__a31o_1
XFILLER_0_152_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12908_ _05655_ _05712_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__xnor2_1
X_19464_ _01297_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__buf_2
X_16676_ _09237_ _09238_ VGND VGND VPWR VPWR _09239_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13888_ _06624_ _06620_ VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__or2_1
XFILLER_0_232_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18415_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[9\] _10364_ _10878_
+ _10879_ _09886_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__o221a_1
X_15627_ _08239_ _08244_ VGND VGND VPWR VPWR _08245_ sky130_fd_sc_hd__or2_1
X_12839_ _05599_ _05600_ _05598_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__o21a_1
X_19395_ _11683_ _11678_ _11696_ _11700_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__nand4_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18346_ _10766_ _10772_ _10811_ VGND VGND VPWR VPWR _10812_ sky130_fd_sc_hd__o21a_1
X_15558_ _08172_ _08177_ _08178_ VGND VGND VPWR VPWR _08180_ sky130_fd_sc_hd__and3_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14509_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[2\] _07078_ _07200_
+ _07201_ VGND VGND VPWR VPWR _07202_ sky130_fd_sc_hd__nand4_2
XFILLER_0_154_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18277_ _10743_ _10744_ VGND VGND VPWR VPWR _10745_ sky130_fd_sc_hd__nor2_1
X_15489_ _08114_ _08128_ VGND VGND VPWR VPWR _08129_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17228_ _09726_ _09758_ VGND VGND VPWR VPWR _09775_ sky130_fd_sc_hd__or2_1
Xinput30 input_tdata[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold803 top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[24\] VGND VGND
+ VPWR VPWR net985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17159_ _09670_ _09680_ _09708_ VGND VGND VPWR VPWR _09709_ sky130_fd_sc_hd__a21o_1
Xhold814 top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[0\] VGND VGND
+ VPWR VPWR net996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 top_inst.axis_in_inst.inbuf_bus\[21\] VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold836 top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[21\] VGND VGND
+ VPWR VPWR net1018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 top_inst.axis_in_inst.inbuf_bus\[16\] VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[11\] VGND VGND
+ VPWR VPWR net1040 sky130_fd_sc_hd__dlygate4sd3_1
X_20170_ _01978_ _01979_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_1000 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold869 top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[25\] VGND VGND
+ VPWR VPWR net1051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_209_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23860_ clknet_leaf_77_clk _00393_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22811_ top_inst.deskew_buff_inst.col_input\[126\] _04476_ _06140_ VGND VGND VPWR
+ VPWR _04478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23791_ clknet_leaf_71_clk _00324_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_211_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22742_ _04268_ _04394_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22673_ _04218_ _04345_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24412_ clknet_leaf_55_clk _00945_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21624_ _03245_ _03353_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__xor2_1
XFILLER_0_164_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24343_ clknet_leaf_8_clk _00876_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[102\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21555_ top_inst.grid_inst.data_path_wires\[17\]\[7\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20506_ _02288_ _02289_ _02241_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__o21a_1
XFILLER_0_160_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21486_ _03176_ _03178_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__and2_1
X_24274_ clknet_leaf_12_clk _00807_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[17\]\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_181_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_244_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23225_ net106 _04714_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__or2_1
X_20437_ _02206_ _02208_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23156_ net485 _04671_ _04681_ _04675_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__o211a_1
X_20368_ _02152_ _02153_ _02154_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__nand3_1
XFILLER_0_28_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22107_ _03770_ _03772_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23087_ net24 _04600_ _04641_ _04632_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20299_ _02086_ _02087_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__xor2_4
XTAP_6346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22038_ _03725_ _03731_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__nand2_1
XTAP_6379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14860_ _07543_ _07542_ VGND VGND VPWR VPWR _07545_ sky130_fd_sc_hd__or2b_1
XTAP_5678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ _06364_ _06553_ VGND VGND VPWR VPWR _06554_ sky130_fd_sc_hd__and2_1
XFILLER_0_230_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14791_ _07446_ _07477_ VGND VGND VPWR VPWR _07478_ sky130_fd_sc_hd__xnor2_2
XTAP_4988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23989_ clknet_leaf_78_clk _00522_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16530_ _09061_ _09062_ _09106_ VGND VGND VPWR VPWR _09107_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_230_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13742_ _06193_ _06214_ _06485_ VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16461_ _09013_ _09012_ VGND VGND VPWR VPWR _09039_ sky130_fd_sc_hd__or2b_1
XFILLER_0_112_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13673_ _06195_ top_inst.grid_inst.data_path_wires\[2\]\[5\] _06210_ _06208_ VGND
+ VGND VPWR VPWR _06419_ sky130_fd_sc_hd__and4_1
XFILLER_0_35_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18200_ _10668_ _10669_ VGND VGND VPWR VPWR _10670_ sky130_fd_sc_hd__xnor2_2
X_15412_ _08053_ _08054_ VGND VGND VPWR VPWR _08055_ sky130_fd_sc_hd__xnor2_1
XPHY_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12624_ _05407_ _05398_ _05435_ _05436_ VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__a211oi_2
X_19180_ _11351_ _11147_ _11520_ _11558_ VGND VGND VPWR VPWR _11597_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16392_ _08959_ _08971_ VGND VGND VPWR VPWR _08972_ sky130_fd_sc_hd__and2b_1
XFILLER_0_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_1279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18131_ _10608_ _10057_ VGND VGND VPWR VPWR _10609_ sky130_fd_sc_hd__or2_1
XPHY_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15343_ _07948_ _07987_ _05335_ VGND VGND VPWR VPWR _07988_ sky130_fd_sc_hd__mux2_1
X_12555_ _05345_ _05369_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__xor2_1
XFILLER_0_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18062_ _10071_ _10561_ _10562_ _10448_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__o211a_1
X_15274_ _07915_ _07919_ VGND VGND VPWR VPWR _07920_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12486_ _05305_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17013_ _09548_ _09565_ _09566_ VGND VGND VPWR VPWR _09567_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14225_ _06932_ _06936_ VGND VGND VPWR VPWR _06937_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14156_ _06825_ _06868_ VGND VGND VPWR VPWR _06870_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_1320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13107_ _05315_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__buf_8
XFILLER_0_238_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14087_ _06801_ _06802_ VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__nor2_1
X_18964_ _11384_ _11385_ VGND VGND VPWR VPWR _11386_ sky130_fd_sc_hd__nand2_1
XFILLER_0_237_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_1416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13038_ _05352_ _05820_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__and2_1
X_17915_ _10035_ _10300_ VGND VGND VPWR VPWR _10420_ sky130_fd_sc_hd__nor2_1
XFILLER_0_225_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18895_ _11273_ _11318_ VGND VGND VPWR VPWR _11319_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17846_ _10327_ _10352_ VGND VGND VPWR VPWR _10353_ sky130_fd_sc_hd__xor2_1
XFILLER_0_206_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_234_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14989_ _07606_ _07627_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _07645_ sky130_fd_sc_hd__and3_1
X_17777_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[9\] _10236_ VGND
+ VGND VPWR VPWR _10285_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19516_ _01347_ _01348_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16728_ _09287_ _09288_ VGND VGND VPWR VPWR _09289_ sky130_fd_sc_hd__nand2_2
XFILLER_0_57_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16659_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[0\] _08183_ _09223_
+ _09184_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__o211a_1
X_19447_ _01268_ _01269_ _01279_ _01280_ VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19378_ _01212_ _01213_ _01214_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18329_ _10790_ _10794_ VGND VGND VPWR VPWR _10795_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_868 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21340_ top_inst.grid_inst.data_path_wires\[17\]\[7\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _03077_ sky130_fd_sc_hd__and3_1
XFILLER_0_167_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21271_ _03008_ _03009_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold600 top_inst.deskew_buff_inst.col_input\[53\] VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[25\] VGND
+ VGND VPWR VPWR net793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold622 top_inst.axis_out_inst.out_buff_data\[78\] VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__dlygate4sd3_1
X_23010_ net616 _04588_ _04597_ _04590_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold633 _00095_ VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__dlygate4sd3_1
X_20222_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _02018_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold644 top_inst.deskew_buff_inst.col_input\[12\] VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold655 top_inst.deskew_buff_inst.col_input\[45\] VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold666 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[2\] VGND
+ VGND VPWR VPWR net848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold677 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[27\] VGND VGND
+ VPWR VPWR net859 sky130_fd_sc_hd__dlygate4sd3_1
X_20153_ _01944_ _01945_ _01963_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__or3b_1
Xhold688 top_inst.axis_out_inst.out_buff_data\[22\] VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[5\] VGND VGND
+ VPWR VPWR net881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20084_ _01896_ _01897_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__xor2_1
XFILLER_0_228_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23912_ clknet_leaf_33_clk _00445_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1083 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23843_ clknet_leaf_96_clk _00376_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23774_ clknet_leaf_63_clk _00307_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20986_ _02725_ _02740_ _02753_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22725_ _04395_ _04396_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_193_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22656_ _04311_ _04330_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21607_ _03336_ _03337_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22587_ _04092_ _04263_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1028 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12340_ _05142_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__clkbuf_2
X_24326_ clknet_leaf_7_clk _00859_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[18\]\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_211_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21538_ _03269_ _03270_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__and2_1
XFILLER_0_209_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24257_ clknet_leaf_110_clk _00790_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_12271_ net698 _05169_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__or2_1
X_21469_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[11\] _03079_ VGND
+ VGND VPWR VPWR _03203_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14010_ _06705_ _06706_ _06726_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23208_ net98 _04701_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__or2_1
X_24188_ clknet_leaf_47_clk _00721_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_31_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23139_ _04658_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__buf_2
XTAP_6121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15961_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[13\] _08452_ VGND
+ VGND VPWR VPWR _08571_ sky130_fd_sc_hd__xnor2_1
XTAP_6165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14912_ _07577_ net229 _07594_ VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__o21a_1
XTAP_5453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17700_ top_inst.grid_inst.data_path_wires\[11\]\[2\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[5\]
+ VGND VGND VPWR VPWR _10210_ sky130_fd_sc_hd__nand2_1
XTAP_5464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15892_ _08451_ _08457_ _08449_ VGND VGND VPWR VPWR _08504_ sky130_fd_sc_hd__a21o_1
X_18680_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[25\] _11116_ net167
+ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__o21a_1
XTAP_5475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14843_ _07241_ _07090_ _07459_ _07496_ VGND VGND VPWR VPWR _07528_ sky130_fd_sc_hd__o211a_1
XTAP_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17631_ _10126_ _10142_ VGND VGND VPWR VPWR _10143_ sky130_fd_sc_hd__xor2_2
XFILLER_0_231_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17562_ _10065_ _10066_ VGND VGND VPWR VPWR _10077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14774_ _07241_ _07242_ _07082_ _07460_ VGND VGND VPWR VPWR _07461_ sky130_fd_sc_hd__or4_4
XFILLER_0_153_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11986_ net820 _05004_ _05006_ _04995_ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_230_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16513_ _09088_ _09089_ VGND VGND VPWR VPWR _09090_ sky130_fd_sc_hd__nand2_1
X_19301_ net193 VGND VGND VPWR VPWR _11700_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13725_ _06465_ _06469_ VGND VGND VPWR VPWR _06470_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_233_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17493_ top_inst.grid_inst.data_path_wires\[11\]\[1\] VGND VGND VPWR VPWR _10025_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_188_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16444_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[11\] _08897_ VGND
+ VGND VPWR VPWR _09023_ sky130_fd_sc_hd__xnor2_1
X_19232_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[15\] _11469_ _11387_
+ VGND VGND VPWR VPWR _11647_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13656_ _06365_ _06360_ _06402_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12607_ _05418_ _05419_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__xnor2_1
X_19163_ _11549_ _11580_ VGND VGND VPWR VPWR _11581_ sky130_fd_sc_hd__xnor2_1
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16375_ _08919_ _08955_ VGND VGND VPWR VPWR _08956_ sky130_fd_sc_hd__xor2_1
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13587_ top_inst.grid_inst.data_path_wires\[2\]\[4\] _06188_ _06210_ _06208_ VGND
+ VGND VPWR VPWR _06335_ sky130_fd_sc_hd__nand4_4
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18114_ _10040_ _10584_ _10596_ _10594_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__o211a_1
X_15326_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[10\] _07924_ _07844_
+ VGND VGND VPWR VPWR _07971_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19094_ _11400_ _11477_ _11438_ VGND VGND VPWR VPWR _11513_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12538_ _05325_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__buf_6
XFILLER_0_186_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18045_ _10545_ _10501_ _10523_ _10530_ VGND VGND VPWR VPWR _10546_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15257_ _07869_ _07903_ VGND VGND VPWR VPWR _07904_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_1138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12469_ _05291_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_151_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14208_ _06919_ _06920_ VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15188_ _07834_ _07835_ VGND VGND VPWR VPWR _07836_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14139_ _06650_ _06628_ VGND VGND VPWR VPWR _06853_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19996_ _01811_ _01812_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_240_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18947_ _11366_ _11369_ VGND VGND VPWR VPWR _11370_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_225_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18878_ top_inst.grid_inst.data_path_wires\[13\]\[6\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[13\]\[7\]
+ VGND VGND VPWR VPWR _11302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17829_ _10037_ _10052_ _10050_ top_inst.grid_inst.data_path_wires\[11\]\[7\] VGND
+ VGND VPWR VPWR _10336_ sky130_fd_sc_hd__a22o_1
XFILLER_0_234_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_233_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20840_ net966 _02491_ _02612_ _02613_ _01863_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__o221a_1
XFILLER_0_77_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20771_ _02516_ _02530_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__or2b_1
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22510_ _04164_ _04167_ _04166_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23490_ clknet_leaf_140_clk net641 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[80\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22441_ _04113_ _04112_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__or2b_1
XFILLER_0_88_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22372_ _04018_ _04017_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__or2b_1
XFILLER_0_72_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24111_ clknet_leaf_16_clk _00644_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_143_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21323_ _03020_ _03022_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24042_ clknet_leaf_42_clk _00575_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21254_ _02964_ _02980_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__nand2_1
Xhold430 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[5\] VGND VGND
+ VPWR VPWR net612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold441 top_inst.axis_out_inst.out_buff_data\[126\] VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold452 _00965_ VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap171 _07180_ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_1
XFILLER_0_25_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold463 top_inst.axis_out_inst.out_buff_data\[73\] VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap182 _06052_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__buf_1
XFILLER_0_64_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20205_ _02004_ _05739_ _02005_ _02006_ VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__o211a_1
Xhold474 _00904_ VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__dlygate4sd3_1
X_21185_ _02924_ _02926_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold485 _00004_ VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[20\] VGND
+ VGND VPWR VPWR net678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20136_ _01932_ _01947_ _05316_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_176_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20067_ _01857_ _01881_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__nand2_1
XTAP_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23826_ clknet_leaf_93_clk _00359_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_11840_ net428 _04912_ _04923_ _04916_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__o211a_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ net364 _04877_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__or2_1
X_23757_ clknet_leaf_135_clk net370 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20969_ _02736_ _02737_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__and2_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[4\] _06242_ _06259_
+ _06260_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__a22o_1
X_22708_ _04354_ _04379_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_971 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _07180_ _07181_ _07182_ VGND VGND VPWR VPWR _07184_ sky130_fd_sc_hd__o21ba_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23688_ clknet_leaf_119_clk _00221_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13441_ _06202_ _05773_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__or2_1
X_22639_ _04306_ _04314_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16160_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[4\] _08745_ VGND
+ VGND VPWR VPWR _08746_ sky130_fd_sc_hd__xor2_2
XFILLER_0_63_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13372_ _06125_ _06127_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__or2b_1
XFILLER_0_51_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15111_ _07758_ _07759_ _07713_ _07715_ VGND VGND VPWR VPWR _07761_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24309_ clknet_leaf_1_clk _00842_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[84\]
+ sky130_fd_sc_hd__dfxtp_1
X_12323_ net926 _05191_ _05199_ _05195_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16091_ _08664_ _08681_ _08687_ _08666_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15042_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[3\] _07673_ _07674_
+ VGND VGND VPWR VPWR _07694_ sky130_fd_sc_hd__a21bo_1
X_12254_ net586 _05156_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19850_ _01652_ _01673_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1060 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12185_ net382 _05115_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18801_ _07707_ VGND VGND VPWR VPWR _11228_ sky130_fd_sc_hd__buf_4
XFILLER_0_222_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19781_ _11703_ _11701_ _11709_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__and3_1
X_16993_ _09545_ _09546_ VGND VGND VPWR VPWR _09547_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18732_ _11164_ _11150_ VGND VGND VPWR VPWR _11165_ sky130_fd_sc_hd__or2_1
XTAP_5250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15944_ _08197_ _08554_ VGND VGND VPWR VPWR _08555_ sky130_fd_sc_hd__and2_1
XTAP_5261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15875_ _08485_ _08486_ VGND VGND VPWR VPWR _08487_ sky130_fd_sc_hd__and2b_1
X_18663_ _10969_ _11102_ _11119_ VGND VGND VPWR VPWR _11120_ sky130_fd_sc_hd__o21a_1
XTAP_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14826_ _07509_ _07510_ _07486_ VGND VGND VPWR VPWR _07512_ sky130_fd_sc_hd__a21oi_1
XTAP_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17614_ _10113_ _10117_ VGND VGND VPWR VPWR _10126_ sky130_fd_sc_hd__and2b_1
XFILLER_0_192_1181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18594_ _11053_ _11016_ VGND VGND VPWR VPWR _11054_ sky130_fd_sc_hd__nand2_1
XTAP_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_231_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14757_ _07400_ _07441_ _07443_ VGND VGND VPWR VPWR _07444_ sky130_fd_sc_hd__a21o_1
X_17545_ _10022_ _10042_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _10062_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_175_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11969_ net849 _04990_ _04997_ _04995_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_137_clk clknet_4_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_137_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_230_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13708_ _06451_ _06452_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__nor2_1
X_17476_ _08870_ _10010_ _10011_ _09231_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14688_ _07328_ _07376_ VGND VGND VPWR VPWR _07377_ sky130_fd_sc_hd__xor2_1
XFILLER_0_184_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19215_ _11594_ _11595_ _11605_ _11603_ VGND VGND VPWR VPWR _11631_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16427_ _08967_ _09005_ VGND VGND VPWR VPWR _09006_ sky130_fd_sc_hd__nor2_2
XFILLER_0_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13639_ _06343_ _06385_ VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16358_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[9\] _08897_ VGND
+ VGND VPWR VPWR _08939_ sky130_fd_sc_hd__xnor2_1
X_19146_ _11522_ _11524_ _11562_ VGND VGND VPWR VPWR _11564_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15309_ _07635_ _07633_ top_inst.grid_inst.data_path_wires\[6\]\[7\] VGND VGND VPWR
+ VPWR _07954_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16289_ _08822_ _08863_ VGND VGND VPWR VPWR _08871_ sky130_fd_sc_hd__nor2_1
X_19077_ _11453_ _11454_ _11496_ VGND VGND VPWR VPWR _11497_ sky130_fd_sc_hd__o21a_1
XFILLER_0_164_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18028_ _10528_ _10529_ VGND VGND VPWR VPWR _10530_ sky130_fd_sc_hd__or2_1
XFILLER_0_199_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19979_ _11177_ _01796_ _01797_ _11714_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22990_ net881 _04583_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__or2_1
XFILLER_0_241_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21941_ _03650_ _03656_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_1038 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21872_ _03566_ _03571_ _03590_ _01984_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__a31o_1
XFILLER_0_210_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23611_ clknet_leaf_104_clk _00144_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20823_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[19\] _02470_ VGND
+ VGND VPWR VPWR _02597_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24591_ clknet_leaf_22_clk _01124_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_33_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_128_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_128_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_171_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23542_ clknet_leaf_129_clk _00075_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20754_ _02516_ _02530_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23473_ clknet_leaf_30_clk net500 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[127\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20685_ _02431_ _02433_ _02430_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22424_ _04025_ _04107_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1036 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22355_ _04038_ _04040_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__xor2_2
XFILLER_0_103_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21306_ _03010_ _03015_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22286_ _03930_ _03931_ _03972_ _06734_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24025_ clknet_4_12__leaf_clk _00558_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold260 _01177_ VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__dlygate4sd3_1
X_21237_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[5\] _02976_ VGND
+ VGND VPWR VPWR _02977_ sky130_fd_sc_hd__xor2_2
Xhold271 _00268_ VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 top_inst.deskew_buff_inst.col_input\[9\] VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold293 _00029_ VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21168_ _02864_ _02885_ _02883_ _02866_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__a22o_1
X_20119_ _01819_ _01930_ _01931_ _01840_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__o211a_1
X_13990_ _06650_ _06618_ VGND VGND VPWR VPWR _06708_ sky130_fd_sc_hd__nand2_1
X_21099_ net1102 _05313_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__nor2_1
X_12941_ _05739_ _05490_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__nand2_1
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15660_ top_inst.grid_inst.data_path_wires\[7\]\[2\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[7\]\[3\]
+ VGND VGND VPWR VPWR _08277_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _05642_ _05671_ _05676_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__nand3_1
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 _05270_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_111 _05313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _07284_ _07301_ VGND VGND VPWR VPWR _07302_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_198_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_122 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23809_ clknet_leaf_74_clk _00342_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11823_ net657 _04903_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__or2_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_clk clknet_4_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _08198_ _08192_ _08210_ VGND VGND VPWR VPWR _08211_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_212_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17330_ _09837_ _09871_ _09836_ VGND VGND VPWR VPWR _09872_ sky130_fd_sc_hd__a21bo_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14542_ _07227_ _07233_ VGND VGND VPWR VPWR _07234_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _04873_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__buf_4
XFILLER_0_139_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _09787_ _09802_ _09803_ _09805_ _09806_ VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__o311a_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _07146_ _07148_ _07165_ _07166_ VGND VGND VPWR VPWR _07167_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16212_ _08764_ _08769_ VGND VGND VPWR VPWR _08796_ sky130_fd_sc_hd__or2b_1
X_19000_ _11420_ _11421_ VGND VGND VPWR VPWR _11422_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13424_ _06190_ _05262_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17192_ _09712_ _09740_ VGND VGND VPWR VPWR _09741_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_1267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16143_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[3\] _08728_ _08729_
+ VGND VGND VPWR VPWR _08730_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13355_ _06100_ _06128_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12306_ net528 _05178_ _05189_ _05182_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__o211a_1
X_16074_ _08673_ _08674_ VGND VGND VPWR VPWR _08675_ sky130_fd_sc_hd__or2_1
X_13286_ _06057_ _06060_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19902_ _01528_ _01722_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__nand2_1
X_15025_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[2\] _07656_ _07657_
+ VGND VGND VPWR VPWR _07678_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_220_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_898 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12237_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[10\] _05143_
+ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19833_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[15\] _01395_ _01396_
+ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__a21o_1
X_12168_ _05044_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_236_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19764_ _01559_ _01591_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16976_ _09529_ _09530_ VGND VGND VPWR VPWR _09531_ sky130_fd_sc_hd__or2_4
X_12099_ _05044_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_194_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18715_ _11152_ _11150_ VGND VGND VPWR VPWR _11153_ sky130_fd_sc_hd__or2_1
Xinput6 input_tdata[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_2
XTAP_5080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15927_ _08530_ _08537_ VGND VGND VPWR VPWR _08538_ sky130_fd_sc_hd__xor2_2
XFILLER_0_223_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19695_ _11684_ _11679_ _11709_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__nand3_4
XFILLER_0_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18646_ _11101_ _11103_ VGND VGND VPWR VPWR _11104_ sky130_fd_sc_hd__xnor2_1
XTAP_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15858_ _08349_ _08393_ _08432_ _08470_ VGND VGND VPWR VPWR _08471_ sky130_fd_sc_hd__a31o_1
X_14809_ _07459_ _07463_ _07461_ VGND VGND VPWR VPWR _07495_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_176_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18577_ _11003_ _10999_ _11036_ _10957_ VGND VGND VPWR VPWR _11038_ sky130_fd_sc_hd__a31o_1
X_15789_ _08354_ _08356_ _08352_ VGND VGND VPWR VPWR _08403_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17528_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _10050_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17459_ _09913_ _09974_ _09994_ VGND VGND VPWR VPWR _09995_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20470_ _02202_ _02225_ _02253_ _02254_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_42_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19129_ _11177_ _11546_ _11547_ _11160_ VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22140_ _03821_ _03830_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__xor2_1
XFILLER_0_113_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22071_ _03762_ _03763_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__xnor2_2
XTAP_6709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21022_ _02786_ _02787_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1096 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_227_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22973_ _04550_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_207_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21924_ _03622_ _03640_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24643_ clknet_leaf_21_clk net609 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[119\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21855_ _03278_ _03573_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20806_ _02517_ _02573_ _02580_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__a21o_1
X_24574_ clknet_leaf_142_clk _01107_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dfxtp_1
X_21786_ _03481_ _03484_ _03505_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_148_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23525_ clknet_leaf_1_clk _00058_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20737_ _02502_ _02504_ VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_203_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23456_ net542 _04840_ _04850_ _04844_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20668_ _02394_ _02414_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22407_ _04089_ _04086_ _04090_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_123_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23387_ net788 _04804_ _04813_ _04808_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20599_ _02352_ _02380_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__xor2_1
X_13140_ net169 _05881_ _05919_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22338_ _03983_ _04023_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__nor2_2
X_13071_ _05851_ _05836_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22269_ _03711_ top_inst.grid_inst.data_path_wires\[18\]\[2\] _03904_ VGND VGND VPWR
+ VPWR _03957_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24008_ clknet_leaf_47_clk _00541_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[9\]
+ sky130_fd_sc_hd__dfxtp_2
X_12022_ net837 _05018_ _05027_ _05022_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16830_ _09369_ _09386_ _09387_ VGND VGND VPWR VPWR _09388_ sky130_fd_sc_hd__nand3_2
XFILLER_0_228_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16761_ _09294_ _09320_ VGND VGND VPWR VPWR _09321_ sky130_fd_sc_hd__xnor2_1
X_13973_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[3\]
+ top_inst.grid_inst.data_path_wires\[3\]\[1\] VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__and3_1
XFILLER_0_219_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18500_ _10948_ _10922_ VGND VGND VPWR VPWR _10962_ sky130_fd_sc_hd__or2b_1
X_12924_ _05701_ _05727_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__xor2_1
X_15712_ _08325_ _08326_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[7\]
+ VGND VGND VPWR VPWR _08328_ sky130_fd_sc_hd__a21oi_1
X_16692_ _09203_ _09187_ _09192_ _09198_ VGND VGND VPWR VPWR _09254_ sky130_fd_sc_hd__a22o_1
X_19480_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _01314_ sky130_fd_sc_hd__inv_2
XFILLER_0_220_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18431_ _10853_ _10894_ VGND VGND VPWR VPWR _10895_ sky130_fd_sc_hd__xor2_1
X_12855_ _05660_ _05661_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__and2_1
XFILLER_0_197_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15643_ _08230_ _08232_ VGND VGND VPWR VPWR _08261_ sky130_fd_sc_hd__or2b_1
XFILLER_0_115_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11806_ net640 _04898_ _04904_ _04902_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15574_ _08180_ _08193_ VGND VGND VPWR VPWR _08195_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18362_ _10741_ _10780_ VGND VGND VPWR VPWR _10828_ sky130_fd_sc_hd__nor2_1
X_12786_ _05327_ _05593_ _05594_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__or3_1
XFILLER_0_139_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17313_ _09726_ _09839_ VGND VGND VPWR VPWR _09856_ sky130_fd_sc_hd__nor2_1
X_14525_ _07215_ _07216_ net171 _07183_ VGND VGND VPWR VPWR _07218_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_138_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _04858_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__buf_8
XFILLER_0_51_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18293_ _10753_ _10759_ VGND VGND VPWR VPWR _10760_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17244_ _09771_ _09773_ VGND VGND VPWR VPWR _09790_ sky130_fd_sc_hd__or2b_1
X_14456_ _07143_ _07144_ _07150_ VGND VGND VPWR VPWR _07151_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13407_ _06170_ _06171_ _06176_ _06178_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17175_ _09625_ _09704_ VGND VGND VPWR VPWR _09724_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14387_ _07087_ _07075_ VGND VGND VPWR VPWR _07088_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16126_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[2\] _08713_ VGND
+ VGND VPWR VPWR _08714_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13338_ _06112_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16057_ _08135_ _06634_ _08662_ _08166_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13269_ _05748_ _05770_ _06043_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15008_ _07655_ _07661_ VGND VGND VPWR VPWR _07662_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19816_ _01629_ _01617_ _01641_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_208_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19747_ _01570_ _01573_ _01574_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__and3_1
X_16959_ _09511_ _09512_ _09510_ VGND VGND VPWR VPWR _09514_ sky130_fd_sc_hd__a21o_1
XFILLER_0_237_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19678_ _01506_ _01507_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__nor2_4
XFILLER_0_116_1008 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18629_ _11076_ _11087_ VGND VGND VPWR VPWR _11088_ sky130_fd_sc_hd__xor2_1
XFILLER_0_177_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21640_ _09787_ _03367_ _03368_ _03369_ _09806_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__o311a_1
XFILLER_0_118_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21571_ _03266_ _03265_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__and2b_1
XANTENNA_11 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_22 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23310_ net537 _04765_ _04770_ _04769_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_33 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20522_ _02224_ _02256_ _02255_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_170_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_44 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24290_ clknet_leaf_120_clk _00823_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_55 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_66 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_244_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_77 net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_209_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23241_ net978 _04726_ _04731_ _04730_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_88 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20453_ _01992_ _02188_ _02237_ _02186_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__a22o_1
XANTENNA_99 _02707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23172_ net870 _04685_ _04692_ _04691_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20384_ _02136_ _02170_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__or2_1
XFILLER_0_207_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22123_ top_inst.grid_inst.data_path_wires\[18\]\[5\] top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[1\]
+ _03697_ top_inst.grid_inst.data_path_wires\[18\]\[6\] VGND VGND VPWR VPWR _03814_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput140 net140 VGND VGND VPWR VPWR output_tdata[77] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput151 net151 VGND VGND VPWR VPWR output_tdata[87] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput162 net162 VGND VGND VPWR VPWR output_tdata[97] sky130_fd_sc_hd__clkbuf_4
XTAP_6528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22054_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[2\] _03726_ _03727_
+ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__a21boi_4
XTAP_6539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21005_ _02718_ _02745_ _02744_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_100_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_242_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22956_ net380 _04557_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21907_ _03611_ _03624_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22887_ net852 _04522_ _04527_ _04524_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_214_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12640_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[5\] _05283_ VGND
+ VGND VPWR VPWR _05452_ sky130_fd_sc_hd__and2_1
X_24626_ clknet_leaf_24_clk net303 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[102\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21838_ _03557_ _03558_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__nor2_1
XFILLER_0_211_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12571_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[0\]
+ _05291_ _05296_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__and4_1
XFILLER_0_148_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24557_ clknet_leaf_135_clk _01090_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dfxtp_4
X_21769_ _03278_ _03492_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__nor2_1
XFILLER_0_194_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_clk clknet_4_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14310_ _07018_ _07019_ VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23508_ clknet_leaf_135_clk net283 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_15290_ _07893_ _07895_ VGND VGND VPWR VPWR _07936_ sky130_fd_sc_hd__or2_1
X_24488_ clknet_leaf_15_clk _01021_ VGND VGND VPWR VPWR top_inst.valid_pipe\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14241_ _06907_ _06952_ VGND VGND VPWR VPWR _06953_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23439_ net711 _04840_ _04841_ _04831_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14172_ _06883_ _06885_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13123_ top_inst.grid_inst.data_path_wires\[1\]\[6\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[1\]\[7\]
+ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18980_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[5\] _11140_ VGND
+ VGND VPWR VPWR _11402_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_237_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _05830_ _05835_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__xnor2_2
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17931_ _10434_ _10410_ VGND VGND VPWR VPWR _10436_ sky130_fd_sc_hd__or2b_1
XFILLER_0_221_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12005_ net862 _05004_ _05017_ _05008_ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__o211a_1
X_17862_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[10\] _10367_ _10283_
+ VGND VGND VPWR VPWR _10368_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19601_ _01426_ _01427_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_219_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16813_ _09198_ _09210_ VGND VGND VPWR VPWR _09371_ sky130_fd_sc_hd__nand2_1
X_17793_ top_inst.grid_inst.data_path_wires\[11\]\[3\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[6\]
+ _10300_ top_inst.grid_inst.data_path_wires\[11\]\[2\] VGND VGND VPWR VPWR _10301_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_156_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_914 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19532_ _01298_ net190 net247 _11703_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__a2bb2o_2
X_16744_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[4\] net1119 net225
+ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _09304_ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13956_ _06671_ _06673_ _06674_ _06675_ VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__and4_1
XFILLER_0_117_1328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12907_ _05709_ _05711_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__xnor2_1
X_19463_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _01297_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16675_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[1\] _09224_ _09225_
+ VGND VGND VPWR VPWR _09238_ sky130_fd_sc_hd__a21boi_1
X_13887_ top_inst.grid_inst.data_path_wires\[3\]\[2\] VGND VGND VPWR VPWR _06624_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18414_ _10835_ _10877_ _09292_ VGND VGND VPWR VPWR _10879_ sky130_fd_sc_hd__a21o_1
X_12838_ _05643_ _05644_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__xnor2_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15626_ _08242_ _08243_ VGND VGND VPWR VPWR _08244_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19394_ _11683_ _11695_ _11700_ _11678_ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__a22o_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18345_ _10726_ _10771_ VGND VGND VPWR VPWR _10811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12769_ _05573_ _05577_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__xor2_1
X_15557_ _08177_ _08178_ _08172_ VGND VGND VPWR VPWR _08179_ sky130_fd_sc_hd__a21oi_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_41_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14508_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[4\] _07068_ _07072_
+ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _07201_ sky130_fd_sc_hd__a22o_1
X_15488_ _08005_ _08104_ _08127_ VGND VGND VPWR VPWR _08128_ sky130_fd_sc_hd__a21oi_1
X_18276_ _10741_ _10742_ _10704_ _10703_ VGND VGND VPWR VPWR _10744_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput20 input_tdata[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
X_17227_ _09771_ _09773_ VGND VGND VPWR VPWR _09774_ sky130_fd_sc_hd__xnor2_2
Xinput31 input_tdata[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_2
X_14439_ _07117_ _07134_ VGND VGND VPWR VPWR _07135_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold804 top_inst.axis_in_inst.inbuf_bus\[29\] VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__dlygate4sd3_1
X_17158_ _09671_ _09679_ VGND VGND VPWR VPWR _09708_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold815 top_inst.deskew_buff_inst.col_input\[59\] VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[13\] VGND VGND
+ VPWR VPWR net1008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold837 top_inst.axis_in_inst.inbuf_bus\[4\] VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold848 top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[28\] VGND VGND
+ VPWR VPWR net1030 sky130_fd_sc_hd__dlygate4sd3_1
X_16109_ _08679_ _08681_ _08699_ _08692_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17089_ _09638_ _09639_ _09635_ VGND VGND VPWR VPWR _09641_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold859 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[0\] VGND VGND
+ VPWR VPWR net1041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_1072 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_244_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22810_ _09787_ _04476_ _04477_ _03929_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23790_ clknet_leaf_70_clk _00323_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_79_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22741_ _04390_ _04411_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_149_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22672_ _04218_ _04345_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24411_ clknet_leaf_55_clk _00944_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21623_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[15\] _03080_ VGND
+ VGND VPWR VPWR _03353_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_clk clknet_4_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24342_ clknet_leaf_8_clk _00875_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[101\]
+ sky130_fd_sc_hd__dfxtp_1
X_21554_ _03284_ _03285_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_776 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20505_ _02003_ top_inst.grid_inst.data_path_wires\[16\]\[6\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[3\]
+ _02051_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__and4_1
X_24273_ clknet_leaf_11_clk _00806_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[17\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21485_ _03210_ _03218_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_133_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_200_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23224_ net763 _04713_ _04721_ _04717_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20436_ _02215_ _02220_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__nor2_1
XFILLER_0_209_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23155_ net74 _04672_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__or2_1
XFILLER_0_219_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20367_ _02109_ _02110_ _02111_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_222_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22106_ _03795_ _03797_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__xnor2_2
XTAP_6314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23086_ net1115 _04602_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_235_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20298_ _02056_ _02059_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__nand2_2
XFILLER_0_100_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_99_clk clknet_4_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22037_ _03725_ _03731_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__or2_1
XTAP_6369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[12\] _06242_ _06551_
+ _06552_ VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__a22o_1
XFILLER_0_242_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14790_ _07475_ _07476_ VGND VGND VPWR VPWR _07477_ sky130_fd_sc_hd__or2_1
XTAP_4978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23988_ clknet_leaf_80_clk _00521_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_230_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13741_ top_inst.grid_inst.data_path_wires\[2\]\[4\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__and2b_1
X_22939_ _04863_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__buf_2
XFILLER_0_230_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16460_ _05440_ _09038_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13672_ _06193_ _06210_ _06208_ _06195_ VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_128_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12623_ _05408_ _05409_ _05434_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__and3_1
X_15411_ _08004_ _08009_ _08007_ VGND VGND VPWR VPWR _08054_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16391_ _08966_ _08970_ VGND VGND VPWR VPWR _08971_ sky130_fd_sc_hd__xor2_1
X_24609_ clknet_leaf_21_clk _01142_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_2_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_23_clk clknet_4_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18130_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _10608_ sky130_fd_sc_hd__clkbuf_4
X_15342_ _07985_ _07986_ VGND VGND VPWR VPWR _07987_ sky130_fd_sc_hd__xnor2_1
XPHY_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12554_ _05362_ _05368_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15273_ _07881_ _07918_ VGND VGND VPWR VPWR _07919_ sky130_fd_sc_hd__xor2_1
X_18061_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[16\] _09494_ VGND
+ VGND VPWR VPWR _10562_ sky130_fd_sc_hd__or2_1
X_12485_ top_inst.skew_buff_inst.row\[0\].output_reg\[7\] top_inst.axis_in_inst.inbuf_bus\[7\]
+ _05267_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__mux2_4
XFILLER_0_48_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17012_ _09562_ _09563_ _09564_ VGND VGND VPWR VPWR _09566_ sky130_fd_sc_hd__a21o_1
X_14224_ net180 _06935_ VGND VGND VPWR VPWR _06936_ sky130_fd_sc_hd__nor2_2
XFILLER_0_145_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14155_ _06825_ _06868_ VGND VGND VPWR VPWR _06869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13106_ _04869_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14086_ _06763_ _06764_ _06762_ VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__o21bai_2
X_18963_ _11336_ _11342_ VGND VGND VPWR VPWR _11385_ sky130_fd_sc_hd__or2b_1
XFILLER_0_120_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13037_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[4\] _05354_ _05818_
+ _05819_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__a22o_1
X_17914_ _10040_ _10054_ VGND VGND VPWR VPWR _10419_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18894_ _11314_ _11317_ VGND VGND VPWR VPWR _11318_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_206_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17845_ _10350_ _10351_ VGND VGND VPWR VPWR _10352_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_238_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17776_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[8\] _10236_ _10283_
+ VGND VGND VPWR VPWR _10284_ sky130_fd_sc_hd__a21o_1
X_14988_ _07624_ _07639_ _07644_ _07643_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19515_ _01299_ _01305_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__or2b_1
X_16727_ _09282_ _09283_ _09286_ VGND VGND VPWR VPWR _09288_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13939_ _05787_ VGND VGND VPWR VPWR _06660_ sky130_fd_sc_hd__buf_4
XFILLER_0_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19446_ _01268_ _01269_ _01279_ _01280_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__nand4_2
X_16658_ _09221_ _09222_ _08181_ VGND VGND VPWR VPWR _09223_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_1303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15609_ _08164_ _08200_ _08227_ VGND VGND VPWR VPWR _08228_ sky130_fd_sc_hd__a21bo_1
X_19377_ _11697_ net243 net191 _11693_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__a22o_1
X_16589_ _09161_ _09162_ VGND VGND VPWR VPWR _09164_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_4_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18328_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[8\] _10793_ VGND
+ VGND VPWR VPWR _10794_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18259_ _10725_ _10726_ VGND VGND VPWR VPWR _10727_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21270_ _02864_ top_inst.grid_inst.data_path_wires\[17\]\[0\] _02895_ _02893_ VGND
+ VGND VPWR VPWR _03009_ sky130_fd_sc_hd__and4_1
XFILLER_0_206_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold601 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[19\] VGND
+ VGND VPWR VPWR net783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold612 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[26\] VGND
+ VGND VPWR VPWR net794 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold623 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[21\] VGND
+ VGND VPWR VPWR net805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20221_ _01997_ _11163_ _02017_ _02006_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold634 top_inst.deskew_buff_inst.col_input\[44\] VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold645 _00211_ VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold656 top_inst.axis_out_inst.out_buff_data\[56\] VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[22\] VGND
+ VGND VPWR VPWR net849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20152_ _01961_ _01962_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__and2_1
Xhold678 top_inst.deskew_buff_inst.col_input\[70\] VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold689 top_inst.deskew_buff_inst.col_input\[40\] VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20083_ _01783_ _01876_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__nor2_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23911_ clknet_leaf_36_clk _00444_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23842_ clknet_leaf_96_clk _00375_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_212_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23773_ clknet_leaf_63_clk _00306_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20985_ _02751_ _02752_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_939 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22724_ _04268_ _04374_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22655_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[21\] _04215_ _04216_
+ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_94_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21606_ _03312_ _03313_ _03335_ VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__nand3_1
XFILLER_0_168_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22586_ _04218_ _04263_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24325_ clknet_leaf_10_clk _00858_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[18\]\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_8_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21537_ _03240_ _03241_ _03268_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__nand3_1
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24256_ clknet_leaf_110_clk _00789_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_12270_ _05142_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__buf_2
X_21468_ _02878_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[2\] _03169_
+ _03168_ _02875_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__a32o_1
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23207_ net845 _04700_ _04711_ _04704_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20419_ _02202_ _02203_ _02185_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24187_ clknet_leaf_47_clk _00720_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_146_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21399_ _02878_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[2\] VGND
+ VGND VPWR VPWR _03135_ sky130_fd_sc_hd__nand2_4
XFILLER_0_31_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23138_ _04655_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23069_ net14 _04628_ _04631_ _04632_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__o211a_1
XTAP_5410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15960_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[12\] _08452_ _08373_
+ VGND VGND VPWR VPWR _08570_ sky130_fd_sc_hd__a21o_1
XTAP_6166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14911_ _05352_ VGND VGND VPWR VPWR _07594_ sky130_fd_sc_hd__buf_2
XTAP_5443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15891_ _08497_ _08502_ VGND VGND VPWR VPWR _08503_ sky130_fd_sc_hd__xnor2_1
XTAP_5476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17630_ _10133_ _10141_ VGND VGND VPWR VPWR _10142_ sky130_fd_sc_hd__xor2_2
X_14842_ _07500_ _07495_ VGND VGND VPWR VPWR _07527_ sky130_fd_sc_hd__and2b_1
XFILLER_0_216_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17561_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[2\] _10075_ VGND
+ VGND VPWR VPWR _10076_ sky130_fd_sc_hd__xor2_1
X_14773_ _07085_ VGND VGND VPWR VPWR _07460_ sky130_fd_sc_hd__inv_2
XFILLER_0_187_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11985_ net730 _04996_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__or2_1
XFILLER_0_231_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19300_ top_inst.skew_buff_inst.row\[3\].output_reg\[5\] top_inst.axis_in_inst.inbuf_bus\[29\]
+ net188 VGND VGND VPWR VPWR _11699_ sky130_fd_sc_hd__mux2_4
XFILLER_0_105_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16512_ _09007_ _09087_ VGND VGND VPWR VPWR _09089_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_230_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13724_ _06467_ _06468_ VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__nor2_1
X_17492_ _10022_ _07611_ _10023_ _10024_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19231_ _11644_ _11597_ VGND VGND VPWR VPWR _11646_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16443_ _08679_ _08688_ _08968_ _08967_ _08677_ VGND VGND VPWR VPWR _09022_ sky130_fd_sc_hd__a32o_1
XFILLER_0_195_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13655_ _06399_ _06401_ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12606_ _05284_ _05292_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__nand2_1
X_19162_ _11578_ _11579_ VGND VGND VPWR VPWR _11580_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16374_ _08920_ _08954_ VGND VGND VPWR VPWR _08955_ sky130_fd_sc_hd__xor2_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13586_ _06188_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[3\]
+ top_inst.grid_inst.data_path_wires\[2\]\[4\] VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__a22o_1
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18113_ _10595_ _08674_ VGND VGND VPWR VPWR _10596_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12537_ _04869_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__buf_8
X_15325_ _07968_ _07969_ VGND VGND VPWR VPWR _07970_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19093_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[11\] _11469_ _11387_
+ VGND VGND VPWR VPWR _11512_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18044_ _10377_ VGND VGND VPWR VPWR _10545_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12468_ top_inst.skew_buff_inst.row\[0\].output_reg\[4\] top_inst.axis_in_inst.inbuf_bus\[4\]
+ net211 VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__mux2_2
X_15256_ _07901_ _07902_ VGND VGND VPWR VPWR _07903_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14207_ _06882_ _06885_ _06881_ VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_151_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15187_ _07622_ _07631_ _07832_ _07833_ VGND VGND VPWR VPWR _07835_ sky130_fd_sc_hd__nand4_4
X_12399_ net346 _05235_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14138_ _06850_ _06851_ VGND VGND VPWR VPWR _06852_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_240_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19995_ _01811_ _01812_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__nor2_2
XFILLER_0_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14069_ top_inst.grid_inst.data_path_wires\[3\]\[7\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _06785_ sky130_fd_sc_hd__and3_1
X_18946_ _11367_ _11368_ VGND VGND VPWR VPWR _11369_ sky130_fd_sc_hd__and2_1
XFILLER_0_225_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18877_ _11276_ _11277_ VGND VGND VPWR VPWR _11301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_241_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17828_ top_inst.grid_inst.data_path_wires\[11\]\[7\] _10052_ _10050_ VGND VGND VPWR
+ VPWR _10335_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17759_ _10059_ _10222_ _10267_ VGND VGND VPWR VPWR _10268_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_162_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20770_ _02508_ _02534_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19429_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[6\] _01262_ _01263_
+ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__and3_1
XFILLER_0_174_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22440_ _03070_ _04122_ _04123_ _03929_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22371_ _04041_ _04015_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__or2b_1
XFILLER_0_45_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24110_ clknet_leaf_14_clk _00643_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_21322_ _03034_ _03059_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24041_ clknet_leaf_42_clk _00574_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold420 top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[1\] VGND VGND
+ VPWR VPWR net602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21253_ _02985_ _02984_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold431 top_inst.axis_out_inst.out_buff_data\[42\] VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold442 top_inst.valid_pipe\[1\] VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold453 top_inst.axis_out_inst.out_buff_data\[117\] VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__dlygate4sd3_1
X_20204_ _10447_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__buf_2
XFILLER_0_102_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap172 _11720_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_1
Xhold464 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[31\] VGND VGND
+ VPWR VPWR net646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold475 top_inst.axis_out_inst.out_buff_data\[88\] VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__dlygate4sd3_1
X_21184_ _02887_ _02925_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__nand2_2
XFILLER_0_141_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold486 top_inst.deskew_buff_inst.col_input\[92\] VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold497 top_inst.axis_out_inst.out_buff_data\[102\] VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20135_ _01924_ _01946_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_244_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20066_ _01879_ _01880_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__and2_1
XTAP_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23825_ clknet_leaf_94_clk _00358_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ net744 _04860_ _04883_ _04875_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__o211a_1
X_23756_ clknet_leaf_135_clk net289 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_20968_ _02715_ _02735_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__nand2_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22707_ _04354_ _04379_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23687_ clknet_leaf_119_clk _00220_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_983 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20899_ _02463_ _02649_ _02503_ VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__a21o_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13440_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _06202_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22638_ _04312_ _04313_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__xor2_1
XFILLER_0_119_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13371_ _06144_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__clkbuf_1
X_22569_ _04225_ _04238_ _04247_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15110_ _07713_ _07715_ _07758_ _07759_ VGND VGND VPWR VPWR _07760_ sky130_fd_sc_hd__a211o_1
X_12322_ net515 _05196_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__or2_1
X_16090_ _08686_ _08684_ VGND VGND VPWR VPWR _08687_ sky130_fd_sc_hd__or2_1
X_24308_ clknet_leaf_2_clk _00841_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[83\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15041_ _07671_ _07692_ VGND VGND VPWR VPWR _07693_ sky130_fd_sc_hd__xor2_2
XFILLER_0_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12253_ net311 _05151_ _05159_ _05155_ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__o211a_1
X_24239_ clknet_leaf_111_clk _00772_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12184_ net350 _05110_ _05119_ _05114_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_1072 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18800_ _11224_ _11225_ _09292_ VGND VGND VPWR VPWR _11227_ sky130_fd_sc_hd__a21o_1
XFILLER_0_236_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19780_ _01534_ _01572_ _01571_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_43_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16992_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[11\] _09419_ VGND
+ VGND VPWR VPWR _09546_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_235_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18731_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _11164_ sky130_fd_sc_hd__buf_2
XFILLER_0_207_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15943_ _08552_ _08553_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[12\]
+ _07816_ VGND VGND VPWR VPWR _08554_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_223_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18662_ _10969_ _11102_ _11101_ VGND VGND VPWR VPWR _11119_ sky130_fd_sc_hd__a21o_1
XTAP_5295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ _08145_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[7\] _08169_
+ top_inst.grid_inst.data_path_wires\[7\]\[5\] VGND VGND VPWR VPWR _08486_ sky130_fd_sc_hd__a22o_1
XTAP_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17613_ _10102_ _10121_ VGND VGND VPWR VPWR _10125_ sky130_fd_sc_hd__nor2_1
X_14825_ _07486_ _07509_ _07510_ VGND VGND VPWR VPWR _07511_ sky130_fd_sc_hd__and3_1
XFILLER_0_215_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18593_ _10595_ _10610_ VGND VGND VPWR VPWR _11053_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ _10022_ _10042_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _10061_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14756_ _07442_ _07398_ _07436_ VGND VGND VPWR VPWR _07443_ sky130_fd_sc_hd__a21oi_1
XTAP_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11968_ net802 _04996_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13707_ top_inst.grid_inst.data_path_wires\[2\]\[4\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[6\]
+ _06450_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17475_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[29\] _09494_ VGND
+ VGND VPWR VPWR _10011_ sky130_fd_sc_hd__or2_1
X_14687_ _07374_ _07375_ VGND VGND VPWR VPWR _07376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11899_ net524 _04951_ _04957_ _04955_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19214_ _11622_ _11629_ VGND VGND VPWR VPWR _11630_ sky130_fd_sc_hd__xor2_2
XFILLER_0_172_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16426_ _08693_ _08690_ _08679_ VGND VGND VPWR VPWR _09005_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_172_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13638_ _06202_ _06200_ top_inst.grid_inst.data_path_wires\[2\]\[7\] VGND VGND VPWR
+ VPWR _06385_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19145_ _11522_ _11524_ _11562_ VGND VGND VPWR VPWR _11563_ sky130_fd_sc_hd__o21ai_1
X_16357_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[8\] _08897_ _08896_
+ VGND VGND VPWR VPWR _08938_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13569_ _06280_ _06279_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15308_ _07915_ _07919_ VGND VGND VPWR VPWR _07953_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19076_ _11455_ _11430_ VGND VGND VPWR VPWR _11496_ sky130_fd_sc_hd__or2b_1
X_16288_ _05732_ VGND VGND VPWR VPWR _08870_ sky130_fd_sc_hd__buf_4
XFILLER_0_112_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18027_ _10283_ _10491_ _10527_ VGND VGND VPWR VPWR _10529_ sky130_fd_sc_hd__nor3_1
XFILLER_0_164_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15239_ _07883_ _07885_ VGND VGND VPWR VPWR _07886_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19978_ net825 _01386_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18929_ _11351_ top_inst.grid_inst.data_path_wires\[13\]\[1\] top_inst.grid_inst.data_path_wires\[13\]\[2\]
+ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[6\] VGND VGND VPWR VPWR
+ _11352_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_226_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_241_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21940_ _03654_ _03655_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__xor2_1
XFILLER_0_171_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21871_ _03566_ _03571_ _03590_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23610_ clknet_leaf_104_clk net446 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20822_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[19\] _02470_ VGND
+ VGND VPWR VPWR _02596_ sky130_fd_sc_hd__nand2_1
X_24590_ clknet_leaf_32_clk _01123_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_72_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23541_ clknet_leaf_128_clk net479 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20753_ _02527_ _02529_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__and2_1
XFILLER_0_175_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23472_ clknet_leaf_32_clk net472 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[126\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20684_ _02462_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__buf_4
XFILLER_0_80_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22423_ _04103_ _04106_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__xor2_1
XFILLER_0_134_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22354_ _03982_ _03998_ _04039_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21305_ _03036_ _03042_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_182_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_206_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22285_ _03930_ _03931_ _03972_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_198_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24024_ clknet_leaf_48_clk _00557_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold250 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[1\] VGND
+ VGND VPWR VPWR net432 sky130_fd_sc_hd__dlygate4sd3_1
X_21236_ _02974_ _02975_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__nand2_1
Xhold261 top_inst.axis_out_inst.out_buff_data\[106\] VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold272 top_inst.deskew_buff_inst.col_input\[64\] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__buf_1
XFILLER_0_178_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold283 _00208_ VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 top_inst.axis_out_inst.out_buff_data\[70\] VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21167_ _02862_ _02887_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_244_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20118_ net756 _01386_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__or2_1
X_21098_ _02850_ _02859_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_176_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12940_ top_inst.grid_inst.data_path_wires\[1\]\[2\] VGND VGND VPWR VPWR _05741_
+ sky130_fd_sc_hd__clkbuf_4
X_20049_ _01834_ _01841_ _01859_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__a21boi_2
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _05642_ _05671_ _05676_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__a21o_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _05275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 _05313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14610_ _07299_ _07300_ VGND VGND VPWR VPWR _07301_ sky130_fd_sc_hd__xor2_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23808_ clknet_leaf_74_clk _00341_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11822_ net865 _04912_ _04913_ _04902_ VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__o211a_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15590_ _08202_ _08209_ VGND VGND VPWR VPWR _08210_ sky130_fd_sc_hd__xnor2_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14541_ _07228_ _07232_ VGND VGND VPWR VPWR _07233_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11753_ _04868_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__buf_6
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23739_ clknet_leaf_127_clk _00272_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17260_ _04869_ VGND VGND VPWR VPWR _09806_ sky130_fd_sc_hd__clkbuf_8
X_14472_ _07163_ _07164_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[5\]
+ VGND VGND VPWR VPWR _07166_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16211_ _08771_ _08777_ VGND VGND VPWR VPWR _08795_ sky130_fd_sc_hd__or2b_1
XFILLER_0_37_975 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13423_ top_inst.grid_inst.data_path_wires\[2\]\[4\] VGND VGND VPWR VPWR _06190_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17191_ _09723_ _09739_ VGND VGND VPWR VPWR _09740_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16142_ _08669_ _08667_ _08686_ _08683_ VGND VGND VPWR VPWR _08729_ sky130_fd_sc_hd__nand4_1
X_13354_ _06125_ _06127_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__xor2_1
XFILLER_0_134_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12305_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[7\] _05183_
+ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13285_ _06057_ _06060_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__nor2_1
X_16073_ _06619_ VGND VGND VPWR VPWR _08674_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19901_ _01528_ _01722_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__nor2_1
X_15024_ _07675_ _07676_ VGND VGND VPWR VPWR _07677_ sky130_fd_sc_hd__or2_1
X_12236_ net464 _05137_ _05149_ _05141_ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19832_ _01611_ _01636_ _01610_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__o21ba_1
X_12167_ net855 _05097_ _05109_ _05101_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19763_ _01560_ _01590_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__xnor2_2
X_16975_ _09527_ _09528_ _09485_ _09487_ VGND VGND VPWR VPWR _09530_ sky130_fd_sc_hd__o211a_1
X_12098_ net538 _05058_ _05070_ _05062_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18714_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _11152_ sky130_fd_sc_hd__clkbuf_4
XTAP_5070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15926_ _08531_ _08536_ VGND VGND VPWR VPWR _08537_ sky130_fd_sc_hd__xnor2_2
X_19694_ _01483_ _01500_ net251 VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__nand3_1
XFILLER_0_127_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 input_tdata[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_4
XTAP_5092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18645_ _10969_ _11102_ VGND VGND VPWR VPWR _11103_ sky130_fd_sc_hd__xor2_1
XTAP_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _08397_ _08391_ _08431_ VGND VGND VPWR VPWR _08470_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_232_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14808_ _07415_ _07465_ VGND VGND VPWR VPWR _07494_ sky130_fd_sc_hd__nand2_1
X_18576_ _11003_ _10999_ _11036_ VGND VGND VPWR VPWR _11037_ sky130_fd_sc_hd__a21oi_1
XTAP_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15788_ _08400_ _08401_ VGND VGND VPWR VPWR _08402_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17527_ _10027_ _10046_ _10048_ _10049_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__o211a_1
X_14739_ _07425_ _07426_ VGND VGND VPWR VPWR _07427_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17458_ _09961_ _09960_ _09976_ VGND VGND VPWR VPWR _09994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16409_ _08986_ _08988_ VGND VGND VPWR VPWR _08989_ sky130_fd_sc_hd__xor2_1
XFILLER_0_145_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17389_ net1051 _09266_ _09927_ _09928_ _09886_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__o221a_1
XFILLER_0_89_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19128_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[12\] _10639_ VGND
+ VGND VPWR VPWR _11547_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19059_ _11400_ _11478_ VGND VGND VPWR VPWR _11479_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_42_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22070_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[3\] _03743_ _03744_
+ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_239_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21021_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[27\] _02468_ VGND
+ VGND VPWR VPWR _02787_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_242_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22972_ top_inst.skew_buff_inst.row\[1\].output_reg\[5\] _04570_ VGND VGND VPWR VPWR
+ _04576_ sky130_fd_sc_hd__or2_1
XFILLER_0_241_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21923_ _03637_ _03639_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24642_ clknet_leaf_30_clk _01175_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[118\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21854_ _03246_ _03573_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__or2_2
XFILLER_0_78_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20805_ _02462_ _02579_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24573_ clknet_leaf_139_clk _01106_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dfxtp_2
X_21785_ net648 _02491_ _03507_ _03508_ _02962_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__o221a_1
XFILLER_0_77_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23524_ clknet_leaf_139_clk net504 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_20736_ net278 _02491_ _02512_ _02513_ _01863_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23455_ top_inst.axis_out_inst.out_buff_data\[115\] _04864_ VGND VGND VPWR VPWR _04850_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_0_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20667_ _02425_ _02446_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__xnor2_1
X_22406_ _04054_ _04085_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_243_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_939 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23386_ net56 _04805_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20598_ _02378_ _02379_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__xnor2_1
X_22337_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[3\]
+ top_inst.grid_inst.data_path_wires\[18\]\[7\] VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13070_ _05829_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__inv_2
X_22268_ _03952_ _03955_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_218_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24007_ clknet_leaf_46_clk _00540_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[8\]
+ sky130_fd_sc_hd__dfxtp_2
X_12021_ net272 _05023_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21219_ _02958_ _02959_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__nor2_1
XFILLER_0_178_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22199_ _03851_ _03855_ _03857_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_79_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16760_ _09318_ _09319_ VGND VGND VPWR VPWR _09320_ sky130_fd_sc_hd__xnor2_2
X_13972_ _06643_ _06624_ VGND VGND VPWR VPWR _06691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_219_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15711_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[7\] _08325_ _08326_
+ VGND VGND VPWR VPWR _08327_ sky130_fd_sc_hd__and3_1
X_12923_ _05656_ _05726_ _05706_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__mux2_1
X_16691_ _09251_ _09252_ VGND VGND VPWR VPWR _09253_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18430_ _10592_ _10892_ _10893_ VGND VGND VPWR VPWR _10894_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_154_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15642_ _08257_ _08259_ VGND VGND VPWR VPWR _08260_ sky130_fd_sc_hd__xnor2_2
X_12854_ _05637_ _05619_ _05659_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__or3_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11805_ top_inst.axis_out_inst.out_buff_data\[80\] _04903_ VGND VGND VPWR VPWR _04904_
+ sky130_fd_sc_hd__or2_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _10825_ _10826_ VGND VGND VPWR VPWR _10827_ sky130_fd_sc_hd__nor2_1
X_15573_ _08180_ _08193_ VGND VGND VPWR VPWR _08194_ sky130_fd_sc_hd__or2_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12785_ _05591_ _05592_ _05556_ _05558_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17312_ _09838_ _09854_ VGND VGND VPWR VPWR _09855_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_138_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14524_ net171 _07183_ _07215_ _07216_ VGND VGND VPWR VPWR _07217_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ top_inst.axis_in_inst.inbuf_valid _04857_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__nand2_8
XFILLER_0_126_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18292_ _10754_ _10758_ VGND VGND VPWR VPWR _10759_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17243_ _09777_ _09780_ VGND VGND VPWR VPWR _09789_ sky130_fd_sc_hd__or2b_1
XFILLER_0_71_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14455_ _07148_ _07149_ VGND VGND VPWR VPWR _07150_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13406_ _05335_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__buf_12
XFILLER_0_148_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17174_ _09701_ _09710_ _09722_ VGND VGND VPWR VPWR _09723_ sky130_fd_sc_hd__a21o_1
XFILLER_0_181_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14386_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _07087_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16125_ _08711_ _08712_ VGND VGND VPWR VPWR _08713_ sky130_fd_sc_hd__nand2_1
X_13337_ _05886_ _06111_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16056_ _08661_ _08140_ VGND VGND VPWR VPWR _08662_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13268_ _05748_ _05770_ _06043_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15007_ _07659_ _07660_ VGND VGND VPWR VPWR _07661_ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12219_ net408 _05137_ _05139_ _05128_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__o211a_1
X_13199_ _05748_ _05765_ _05763_ _05750_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_196_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19815_ _01631_ _01640_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16958_ _09510_ _09511_ _09512_ VGND VGND VPWR VPWR _09513_ sky130_fd_sc_hd__nand3_1
X_19746_ _01571_ _01572_ _01534_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__a21o_1
XFILLER_0_223_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15909_ _08149_ _08169_ _08518_ VGND VGND VPWR VPWR _08520_ sky130_fd_sc_hd__a21oi_1
X_19677_ _01504_ _01505_ _01476_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__a21oi_1
X_16889_ _09413_ _09445_ VGND VGND VPWR VPWR _09446_ sky130_fd_sc_hd__xor2_1
XFILLER_0_204_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18628_ _11085_ _11086_ VGND VGND VPWR VPWR _11087_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18559_ _11018_ _11019_ VGND VGND VPWR VPWR _11020_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21570_ _03280_ _03301_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_12 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_23 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20521_ _02303_ _02304_ VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__nor2_1
XANTENNA_34 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_45 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_67 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23240_ net113 _04727_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_78 net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20452_ _01992_ _02020_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_89 net139 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23171_ net80 _04687_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20383_ _02168_ _02169_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__xor2_1
XFILLER_0_141_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22122_ _03780_ _03783_ _03782_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput130 net130 VGND VGND VPWR VPWR output_tdata[68] sky130_fd_sc_hd__clkbuf_4
Xoutput141 net141 VGND VGND VPWR VPWR output_tdata[78] sky130_fd_sc_hd__clkbuf_4
Xoutput152 net152 VGND VGND VPWR VPWR output_tdata[88] sky130_fd_sc_hd__clkbuf_4
XTAP_6507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput163 net163 VGND VGND VPWR VPWR output_tdata[98] sky130_fd_sc_hd__clkbuf_4
XTAP_6518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22053_ _03745_ _03746_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__or2_2
XTAP_6529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21004_ _02769_ _02770_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_220_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_216_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22955_ net612 _04562_ _04566_ _04564_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_242_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21906_ _03622_ _03623_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22886_ top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[0\] _04517_ VGND
+ VGND VPWR VPWR _04527_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24625_ clknet_leaf_25_clk net425 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[101\]
+ sky130_fd_sc_hd__dfxtp_1
X_21837_ _03279_ _03556_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12570_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[2\] _05283_ _05364_
+ _05363_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__a31o_1
X_24556_ clknet_leaf_136_clk _01089_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dfxtp_2
X_21768_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[21\] _03122_ VGND
+ VGND VPWR VPWR _03492_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23507_ clknet_leaf_136_clk net326 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20719_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[15\] _02470_ VGND
+ VGND VPWR VPWR _02497_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24487_ clknet_leaf_84_clk _01020_ VGND VGND VPWR VPWR top_inst.valid_pipe\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21699_ _03278_ _03424_ VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14240_ _06950_ _06951_ VGND VGND VPWR VPWR _06952_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23438_ net444 _04835_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14171_ _06842_ _06844_ _06884_ VGND VGND VPWR VPWR _06885_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_151_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23369_ net48 _04792_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13122_ _05858_ _05860_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13053_ _05831_ _05834_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__xor2_2
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17930_ _10410_ _10434_ VGND VGND VPWR VPWR _10435_ sky130_fd_sc_hd__or2b_1
XFILLER_0_30_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12004_ net458 _05010_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__or2_1
X_17861_ _10236_ VGND VGND VPWR VPWR _10367_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_187_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16812_ _09335_ _09336_ _09339_ VGND VGND VPWR VPWR _09370_ sky130_fd_sc_hd__and3_1
X_19600_ _11177_ _01430_ _01431_ _11714_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17792_ _10059_ VGND VGND VPWR VPWR _10300_ sky130_fd_sc_hd__inv_2
XFILLER_0_219_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_205_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19531_ _01297_ _01314_ _11681_ net246 VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__or4b_4
X_16743_ _09300_ _09301_ _09295_ VGND VGND VPWR VPWR _09303_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13955_ _06661_ _06672_ VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__or2_1
XFILLER_0_221_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12906_ _05658_ _05684_ _05710_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__o21ai_1
X_19462_ _01296_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16674_ _09235_ _09236_ VGND VGND VPWR VPWR _09237_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13886_ _06184_ _06192_ _06623_ _06446_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18413_ _10835_ _10877_ VGND VGND VPWR VPWR _10878_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15625_ _08143_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[2\] _08240_
+ _08241_ VGND VGND VPWR VPWR _08243_ sky130_fd_sc_hd__nand4_2
X_12837_ _05298_ _05306_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__nand2_2
X_19393_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[4\] _01203_ _01204_
+ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_9_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18344_ _10801_ _10809_ VGND VGND VPWR VPWR _10810_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_201_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15556_ _08175_ _08176_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[1\]
+ VGND VGND VPWR VPWR _08178_ sky130_fd_sc_hd__a21o_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _05538_ _05576_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[3\]
+ _07068_ _07072_ VGND VGND VPWR VPWR _07200_ sky130_fd_sc_hd__nand4_2
XFILLER_0_173_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18275_ _10704_ _10703_ _10741_ _10742_ VGND VGND VPWR VPWR _10743_ sky130_fd_sc_hd__and4bb_1
X_15487_ _08005_ _08104_ _08103_ VGND VGND VPWR VPWR _08127_ sky130_fd_sc_hd__o21a_1
X_12699_ _05507_ _05508_ _05506_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17226_ _09624_ _09772_ VGND VGND VPWR VPWR _09773_ sky130_fd_sc_hd__xor2_2
XFILLER_0_116_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14438_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[3\] _07133_ _06701_
+ VGND VGND VPWR VPWR _07134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput10 input_tdata[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_4
Xinput21 input_tdata[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_25_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput32 input_tdata[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17157_ _09702_ _09706_ VGND VGND VPWR VPWR _09707_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold805 top_inst.axis_in_inst.inbuf_bus\[24\] VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__dlygate4sd3_1
X_14369_ _07072_ VGND VGND VPWR VPWR _07073_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold816 top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[14\] VGND VGND
+ VPWR VPWR net998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16108_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[7\] _08684_ VGND
+ VGND VPWR VPWR _08699_ sky130_fd_sc_hd__or2_1
Xhold827 top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[23\] VGND VGND
+ VPWR VPWR net1009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 _00978_ VGND VGND VPWR VPWR net1020 sky130_fd_sc_hd__dlygate4sd3_1
X_17088_ _09635_ _09638_ _09639_ VGND VGND VPWR VPWR _09640_ sky130_fd_sc_hd__and3_1
Xhold849 top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[3\] VGND VGND
+ VPWR VPWR net1031 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16039_ _08620_ _08621_ _08646_ _08618_ VGND VGND VPWR VPWR _08647_ sky130_fd_sc_hd__a211o_1
XFILLER_0_161_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_224_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_237_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19729_ net826 _01386_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__or2_1
XFILLER_0_237_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22740_ _04410_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22671_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[23\] _04163_ VGND
+ VGND VPWR VPWR _04345_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24410_ clknet_leaf_57_clk _00943_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21622_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[14\] _03122_ _03123_
+ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24341_ clknet_leaf_8_clk _00874_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[100\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21553_ _03281_ _03283_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20504_ top_inst.grid_inst.data_path_wires\[16\]\[6\] _02013_ _02011_ _02003_ VGND
+ VGND VPWR VPWR _02288_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_133_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24272_ clknet_leaf_97_clk _00805_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21484_ _03215_ _03217_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__xor2_2
XFILLER_0_105_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23223_ net105 _04714_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20435_ _02168_ _02175_ _02170_ _02136_ _02216_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__o221a_1
XFILLER_0_209_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23154_ net832 _04671_ _04680_ _04675_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__o211a_1
X_20366_ _02150_ _02151_ _02149_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__a21o_1
XFILLER_0_219_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22105_ _03762_ _03763_ _03796_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__a21o_1
XTAP_6304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23085_ net22 _04628_ _04640_ _04632_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__o211a_1
X_20297_ _02076_ _02085_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__xnor2_4
XTAP_6326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22036_ _03729_ _03730_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__xnor2_1
XTAP_6359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23987_ clknet_leaf_80_clk _00520_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_199_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13740_ _06477_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__inv_2
XFILLER_0_225_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22938_ net1037 _04548_ _04556_ _04551_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13671_ _06415_ _06416_ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__xor2_1
XFILLER_0_211_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22869_ _06619_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__buf_2
XFILLER_0_116_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15410_ _08051_ _08052_ VGND VGND VPWR VPWR _08053_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12622_ _05408_ _05409_ _05434_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__a21oi_2
X_24608_ clknet_leaf_22_clk _01141_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_38_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16390_ _08932_ _08969_ VGND VGND VPWR VPWR _08970_ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15341_ _07941_ _07943_ _07939_ VGND VGND VPWR VPWR _07986_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12553_ _05365_ _05367_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__nor2_1
X_24539_ clknet_leaf_130_clk _01072_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_87_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18060_ _10544_ _10560_ VGND VGND VPWR VPWR _10561_ sky130_fd_sc_hd__xor2_1
X_15272_ _07622_ _07916_ _07917_ VGND VGND VPWR VPWR _07918_ sky130_fd_sc_hd__a21bo_1
X_12484_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _05304_ sky130_fd_sc_hd__buf_2
X_17011_ _09562_ _09563_ _09564_ VGND VGND VPWR VPWR _09565_ sky130_fd_sc_hd__nand3_2
XFILLER_0_22_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14223_ _06898_ _06933_ _06860_ VGND VGND VPWR VPWR _06935_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14154_ _06867_ _06818_ VGND VGND VPWR VPWR _06868_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13105_ _05885_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_238_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14085_ _06798_ _06800_ VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__xnor2_2
X_18962_ _11341_ _11337_ VGND VGND VPWR VPWR _11384_ sky130_fd_sc_hd__or2b_1
XFILLER_0_24_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13036_ _05800_ _05817_ _05315_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__o21a_1
X_17913_ _10411_ _10417_ VGND VGND VPWR VPWR _10418_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_237_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18893_ _11315_ _11316_ VGND VGND VPWR VPWR _11317_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_206_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17844_ _10289_ _10309_ _10307_ VGND VGND VPWR VPWR _10351_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_206_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17775_ _10235_ VGND VGND VPWR VPWR _10283_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_234_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14987_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[7\] _07641_ VGND
+ VGND VPWR VPWR _07644_ sky130_fd_sc_hd__or2_1
XFILLER_0_206_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16726_ _09282_ _09283_ _09286_ VGND VGND VPWR VPWR _09287_ sky130_fd_sc_hd__nand3_2
X_19514_ _01304_ _01300_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__or2b_1
X_13938_ _06658_ _06659_ _05440_ VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19445_ _01277_ _01278_ _01242_ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16657_ _09189_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[0\] _09187_
+ VGND VGND VPWR VPWR _09222_ sky130_fd_sc_hd__and3_1
XFILLER_0_187_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13869_ _06540_ _06602_ _06605_ VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__and3_1
XFILLER_0_201_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15608_ top_inst.grid_inst.data_path_wires\[7\]\[0\] _08164_ _08161_ top_inst.grid_inst.data_path_wires\[7\]\[1\]
+ VGND VGND VPWR VPWR _08227_ sky130_fd_sc_hd__a22o_1
X_19376_ _11697_ _11693_ net243 net191 VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__nand4_2
XFILLER_0_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16588_ _09161_ _09162_ VGND VGND VPWR VPWR _09163_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18327_ _10791_ _10792_ VGND VGND VPWR VPWR _10793_ sky130_fd_sc_hd__nor2_4
X_15539_ _07617_ VGND VGND VPWR VPWR _08166_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18258_ _10599_ top_inst.grid_inst.data_path_wires\[12\]\[0\] _10612_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[5\]
+ VGND VGND VPWR VPWR _10726_ sky130_fd_sc_hd__and4_2
XFILLER_0_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17209_ _09755_ _09756_ VGND VGND VPWR VPWR _09757_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18189_ _10657_ _10658_ _10642_ VGND VGND VPWR VPWR _10660_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold602 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[4\] VGND VGND
+ VPWR VPWR net784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold613 top_inst.deskew_buff_inst.col_input\[43\] VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__dlygate4sd3_1
X_20220_ _02016_ _11689_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold624 _00092_ VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 top_inst.deskew_buff_inst.col_input\[104\] VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold646 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[5\] VGND VGND
+ VPWR VPWR net828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 top_inst.deskew_buff_inst.col_input\[76\] VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[7\] VGND VGND
+ VPWR VPWR net850 sky130_fd_sc_hd__dlygate4sd3_1
X_20151_ _01959_ _01960_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold679 top_inst.deskew_buff_inst.col_input\[52\] VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20082_ _01891_ _01895_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__xor2_4
XFILLER_0_176_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23910_ clknet_leaf_36_clk _00443_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23841_ clknet_leaf_96_clk _00374_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_240_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23772_ clknet_leaf_63_clk _00305_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_20984_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[23\] _02559_ _02722_
+ _02720_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__a31o_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22723_ _04394_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__inv_2
XFILLER_0_220_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22654_ _04307_ _04310_ _04309_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_34_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21605_ _03312_ _03313_ _03335_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__a21o_1
XFILLER_0_192_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22585_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[19\] _04163_ VGND
+ VGND VPWR VPWR _04263_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24324_ clknet_leaf_10_clk _00857_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[18\]\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_168_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21536_ _03240_ _03241_ _03268_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24255_ clknet_leaf_110_clk _00788_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_21467_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[10\] _03080_ _03123_
+ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__a21o_1
XFILLER_0_209_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23206_ net97 _04701_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__or2_1
X_20418_ _02185_ _02202_ _02203_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24186_ clknet_leaf_47_clk _00719_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_21398_ _03131_ _03133_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23137_ net661 _04656_ _04670_ _04662_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__o211a_1
X_20349_ _02066_ _02128_ _02127_ _02131_ _02099_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_219_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23068_ _04550_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__clkbuf_4
XTAP_5400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14910_ _07592_ VGND VGND VPWR VPWR _07593_ sky130_fd_sc_hd__buf_6
XTAP_5433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22019_ _03698_ _03680_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__a21oi_1
XTAP_6189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15890_ _08498_ _08501_ VGND VGND VPWR VPWR _08502_ sky130_fd_sc_hd__xor2_1
XTAP_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ _07521_ _07525_ VGND VGND VPWR VPWR _07526_ sky130_fd_sc_hd__xnor2_1
XTAP_5488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ _10073_ _10074_ VGND VGND VPWR VPWR _10075_ sky130_fd_sc_hd__nand2_1
X_14772_ _07083_ _07090_ VGND VGND VPWR VPWR _07459_ sky130_fd_sc_hd__nand2_2
XTAP_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11984_ net598 _05004_ _05005_ _04995_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__o211a_1
XFILLER_0_230_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16511_ _09007_ _09087_ VGND VGND VPWR VPWR _09088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13723_ _06385_ _06466_ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__and2_1
X_17491_ _07617_ VGND VGND VPWR VPWR _10024_ sky130_fd_sc_hd__buf_2
XFILLER_0_105_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19230_ _11644_ _11600_ _11622_ _11629_ VGND VGND VPWR VPWR _11645_ sky130_fd_sc_hd__o2bb2a_1
X_16442_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[10\] _08975_ _08896_
+ VGND VGND VPWR VPWR _09021_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13654_ _06350_ _06352_ _06400_ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_73_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12605_ _05416_ _05417_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__nor2_1
X_19161_ _11576_ _11577_ VGND VGND VPWR VPWR _11579_ sky130_fd_sc_hd__nand2_1
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16373_ _08952_ _08953_ VGND VGND VPWR VPWR _08954_ sky130_fd_sc_hd__or2_1
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13585_ _06296_ _06332_ VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__xor2_1
XFILLER_0_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18112_ top_inst.grid_inst.data_path_wires\[12\]\[7\] VGND VGND VPWR VPWR _10595_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15324_ _07952_ _07953_ _07967_ VGND VGND VPWR VPWR _07969_ sky130_fd_sc_hd__nand3_1
X_12536_ net1048 _05314_ _05351_ _05308_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19092_ _11476_ _11491_ _11510_ VGND VGND VPWR VPWR _11511_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_124_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18043_ _10486_ _10516_ _10539_ _10543_ _10538_ VGND VGND VPWR VPWR _10544_ sky130_fd_sc_hd__a32o_1
X_15255_ _07898_ _07900_ VGND VGND VPWR VPWR _07902_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12467_ _05269_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14206_ _06917_ _06918_ VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15186_ _07621_ _07631_ _07832_ _07833_ VGND VGND VPWR VPWR _07834_ sky130_fd_sc_hd__a22o_1
X_12398_ net505 _05230_ _05241_ _05234_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__o211a_1
XFILLER_0_238_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14137_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[3\]\[3\]
+ _06849_ VGND VGND VPWR VPWR _06851_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19994_ _01778_ _01785_ _01807_ _01769_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_240_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_1327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14068_ top_inst.grid_inst.data_path_wires\[3\]\[6\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[3\]\[7\]
+ VGND VGND VPWR VPWR _06784_ sky130_fd_sc_hd__a22o_1
X_18945_ _11323_ _11298_ VGND VGND VPWR VPWR _11368_ sky130_fd_sc_hd__or2b_1
XFILLER_0_238_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13019_ _05791_ _05796_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18876_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[6\] _11265_ _11266_
+ VGND VGND VPWR VPWR _11300_ sky130_fd_sc_hd__a21bo_1
XTAP_6690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17827_ _10297_ _10305_ VGND VGND VPWR VPWR _10334_ sky130_fd_sc_hd__or2b_1
XFILLER_0_233_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17758_ _10221_ _10220_ VGND VGND VPWR VPWR _10267_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16709_ _09267_ _09268_ _09269_ VGND VGND VPWR VPWR _09270_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_89_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17689_ top_inst.grid_inst.data_path_wires\[11\]\[7\] _10037_ _10044_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _10199_ sky130_fd_sc_hd__nand4_1
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19428_ _11683_ _11678_ _11700_ _11705_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__nand4_1
XFILLER_0_134_1281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19359_ _01178_ _01195_ _01196_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22370_ _04040_ _04038_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__or2b_1
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21321_ _03035_ _03058_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24040_ clknet_leaf_42_clk _00573_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold410 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[11\] VGND
+ VGND VPWR VPWR net592 sky130_fd_sc_hd__dlygate4sd3_1
X_21252_ _02991_ VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold421 _00959_ VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[15\] VGND
+ VGND VPWR VPWR net614 sky130_fd_sc_hd__dlygate4sd3_1
X_20203_ _04858_ _11709_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__or2_2
Xhold443 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[0\] VGND
+ VGND VPWR VPWR net625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 top_inst.deskew_buff_inst.col_input\[86\] VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap173 _07101_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__buf_1
XFILLER_0_13_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21183_ top_inst.grid_inst.data_path_wires\[17\]\[1\] top_inst.grid_inst.data_path_wires\[17\]\[0\]
+ _02889_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__and3_1
Xhold465 top_inst.deskew_buff_inst.col_input\[55\] VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold476 top_inst.axis_out_inst.out_buff_data\[86\] VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _00067_ VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20134_ _01944_ _01945_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__xor2_1
Xhold498 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[28\] VGND
+ VGND VPWR VPWR net680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20065_ _01853_ _01878_ _01869_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__nand3_1
XFILLER_0_77_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23824_ clknet_leaf_94_clk _00357_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23755_ clknet_leaf_135_clk net277 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20967_ _02715_ _02735_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__or2_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22706_ _04377_ _04378_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23686_ clknet_leaf_118_clk _00219_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20898_ _02518_ _02668_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22637_ _04137_ _04293_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13370_ _05886_ _06143_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__and2_1
X_22568_ _04239_ _04246_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_228_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24307_ clknet_leaf_2_clk _00840_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[82\]
+ sky130_fd_sc_hd__dfxtp_1
X_12321_ net824 _05191_ _05198_ _05195_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21519_ top_inst.grid_inst.data_path_wires\[17\]\[7\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[5\]
+ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22499_ _04160_ _04156_ _04180_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__a21oi_1
X_15040_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[4\] _07691_ VGND
+ VGND VPWR VPWR _07692_ sky130_fd_sc_hd__xor2_2
X_12252_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[16\] _05156_
+ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__or2_1
X_24238_ clknet_leaf_111_clk _00771_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12183_ top_inst.axis_out_inst.out_buff_data\[19\] _05115_ VGND VGND VPWR VPWR _05119_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_82_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24169_ clknet_leaf_23_clk _00702_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16991_ _09198_ _09219_ _09507_ _09506_ _09207_ VGND VGND VPWR VPWR _09545_ sky130_fd_sc_hd__a32o_1
XFILLER_0_236_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18730_ _05755_ VGND VGND VPWR VPWR _11163_ sky130_fd_sc_hd__buf_4
X_15942_ _08549_ _08551_ _06404_ VGND VGND VPWR VPWR _08553_ sky130_fd_sc_hd__a21o_1
XTAP_5230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18661_ _11099_ _11105_ _11107_ VGND VGND VPWR VPWR _11118_ sky130_fd_sc_hd__o21a_1
XFILLER_0_235_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ top_inst.grid_inst.data_path_wires\[7\]\[5\] _08145_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[7\]
+ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[6\] VGND VGND VPWR VPWR
+ _08485_ sky130_fd_sc_hd__and4_1
XFILLER_0_244_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14824_ _07467_ _07470_ _07508_ VGND VGND VPWR VPWR _07510_ sky130_fd_sc_hd__nand3_1
XTAP_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17612_ net1053 _09266_ _10123_ _10124_ _09886_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__o221a_1
XTAP_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18592_ _10595_ _10857_ _10975_ _11013_ VGND VGND VPWR VPWR _11052_ sky130_fd_sc_hd__o211a_1
XTAP_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_230_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17543_ _10040_ _10046_ _10060_ _10049_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14755_ _07361_ _07362_ _07394_ _07395_ VGND VGND VPWR VPWR _07442_ sky130_fd_sc_hd__a211o_1
XTAP_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ _04876_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__buf_2
XFILLER_0_54_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13706_ _06190_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[6\] _06450_
+ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17474_ _09990_ _10000_ _10008_ _10009_ VGND VGND VPWR VPWR _10010_ sky130_fd_sc_hd__and4_1
X_14686_ _07079_ _07074_ _07086_ _07090_ VGND VGND VPWR VPWR _07375_ sky130_fd_sc_hd__nand4_1
XFILLER_0_54_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11898_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[24\] _04956_
+ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16425_ _08966_ _08970_ VGND VGND VPWR VPWR _09004_ sky130_fd_sc_hd__nand2_1
X_19213_ _11627_ _11628_ VGND VGND VPWR VPWR _11629_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13637_ _06196_ _06343_ VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19144_ _11520_ _11561_ VGND VGND VPWR VPWR _11562_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16356_ _08934_ _08936_ VGND VGND VPWR VPWR _08937_ sky130_fd_sc_hd__xnor2_1
X_13568_ _06278_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15307_ _07914_ _07913_ VGND VGND VPWR VPWR _07952_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12519_ _05335_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__buf_4
X_19075_ _11468_ _11494_ VGND VGND VPWR VPWR _11495_ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16287_ _08869_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13499_ _06244_ _06249_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18026_ _10283_ _10491_ _10527_ VGND VGND VPWR VPWR _10528_ sky130_fd_sc_hd__o21a_1
XFILLER_0_242_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15238_ _07831_ _07834_ _07835_ _07884_ _07828_ VGND VGND VPWR VPWR _07885_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15169_ _07117_ _07817_ VGND VGND VPWR VPWR _07818_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19977_ _01792_ _01795_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__xor2_2
XFILLER_0_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18928_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _11351_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18859_ _11262_ _11282_ _11283_ VGND VGND VPWR VPWR _11284_ sky130_fd_sc_hd__and3_1
XFILLER_0_179_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21870_ _03563_ _03589_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20821_ _02463_ _02579_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23540_ clknet_leaf_128_clk net482 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20752_ _02528_ _02519_ _02526_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__nand3_1
XFILLER_0_72_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23471_ clknet_leaf_31_clk net667 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[125\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20683_ _02460_ _02461_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22422_ _04104_ _04070_ _04105_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_190_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22353_ _03995_ _03997_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21304_ _03037_ _03041_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__xor2_2
X_22284_ _03932_ _03971_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24023_ clknet_leaf_53_clk _00556_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21235_ _02873_ top_inst.grid_inst.data_path_wires\[17\]\[4\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[1\]
+ _02882_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__nand4_1
Xhold240 top_inst.axis_out_inst.out_buff_data\[4\] VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 _00168_ VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 top_inst.axis_out_inst.out_buff_data\[107\] VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold273 _00039_ VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21166_ net325 _06169_ _02908_ _02909_ VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__o211a_1
Xhold284 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[1\] VGND
+ VGND VPWR VPWR net466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 top_inst.deskew_buff_inst.col_input\[58\] VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20117_ _01912_ _01929_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__xor2_2
XFILLER_0_244_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1055 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21097_ _02857_ _02858_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_244_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20048_ net1099 _01202_ _01861_ _01862_ _01863_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__o221a_1
XFILLER_0_137_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12870_ _05644_ _05675_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _05275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_113 _05313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23807_ clknet_leaf_74_clk _00340_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11821_ net629 _04903_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__or2_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21999_ _03682_ _02881_ _03701_ _03702_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14540_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[7\] _07231_ VGND
+ VGND VPWR VPWR _07232_ sky130_fd_sc_hd__xor2_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11752_ net410 _04865_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23738_ clknet_leaf_127_clk net569 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_230_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[5\] _07163_ _07164_
+ VGND VGND VPWR VPWR _07165_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23669_ clknet_leaf_116_clk net344 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16210_ _08776_ _08772_ VGND VGND VPWR VPWR _08794_ sky130_fd_sc_hd__or2b_1
XFILLER_0_138_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13422_ _05744_ _05256_ _06189_ _06183_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__o211a_1
X_17190_ _09725_ _09738_ VGND VGND VPWR VPWR _09739_ sky130_fd_sc_hd__xor2_1
XFILLER_0_153_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16141_ _08667_ _08686_ _08683_ _08669_ VGND VGND VPWR VPWR _08728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13353_ _06054_ _06091_ _06126_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12304_ net554 _05178_ _05188_ _05182_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16072_ top_inst.grid_inst.data_path_wires\[8\]\[5\] VGND VGND VPWR VPWR _08673_
+ sky130_fd_sc_hd__clkbuf_4
X_13284_ _06058_ _06019_ _06059_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19900_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[19\] _01480_ VGND
+ VGND VPWR VPWR _01722_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_161_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15023_ _07673_ _07674_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[3\]
+ VGND VGND VPWR VPWR _07676_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12235_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[9\] _05143_
+ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__or2_1
X_19831_ _01633_ _01635_ _01655_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__a21o_1
XFILLER_0_236_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12166_ net618 _05102_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__or2_1
XFILLER_0_235_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19762_ _01588_ _01589_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__xor2_2
X_16974_ _09485_ _09487_ _09527_ _09528_ VGND VGND VPWR VPWR _09529_ sky130_fd_sc_hd__a211oi_2
X_12097_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[14\] _05063_
+ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__or2_1
XFILLER_0_159_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18713_ _11130_ _10607_ _11151_ _11137_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__o211a_1
XTAP_5060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15925_ _08534_ _08535_ VGND VGND VPWR VPWR _08536_ sky130_fd_sc_hd__nor2_1
XFILLER_0_223_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19693_ _01478_ _01482_ _01521_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__a21o_1
Xinput8 input_tdata[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XTAP_5082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15856_ _08467_ _08468_ VGND VGND VPWR VPWR _08469_ sky130_fd_sc_hd__nor2_1
X_18644_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[16\] _10923_ VGND
+ VGND VPWR VPWR _11102_ sky130_fd_sc_hd__xnor2_2
XTAP_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14807_ _07464_ _07458_ VGND VGND VPWR VPWR _07493_ sky130_fd_sc_hd__or2b_1
XFILLER_0_59_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_231_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15787_ _08163_ _08167_ VGND VGND VPWR VPWR _08401_ sky130_fd_sc_hd__nand2_1
X_18575_ _11004_ _11035_ VGND VGND VPWR VPWR _11036_ sky130_fd_sc_hd__xnor2_1
X_12999_ _05734_ _05761_ _05783_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__a21oi_1
XTAP_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14738_ _07410_ _07411_ _07424_ VGND VGND VPWR VPWR _07426_ sky130_fd_sc_hd__nand3_1
XFILLER_0_146_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17526_ _07617_ VGND VGND VPWR VPWR _10049_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17457_ _09919_ _09957_ _09976_ VGND VGND VPWR VPWR _09993_ sky130_fd_sc_hd__and3b_1
XFILLER_0_184_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14669_ _07308_ _07309_ _07354_ VGND VGND VPWR VPWR _07358_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16408_ _08947_ _08948_ _08987_ VGND VGND VPWR VPWR _08988_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17388_ _09908_ _09909_ _09926_ _07439_ VGND VGND VPWR VPWR _09928_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16339_ _08910_ _08912_ VGND VGND VPWR VPWR _08920_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19127_ _11544_ _11545_ VGND VGND VPWR VPWR _11546_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19058_ _11438_ _11477_ VGND VGND VPWR VPWR _11478_ sky130_fd_sc_hd__nor2_2
XFILLER_0_140_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18009_ _10475_ VGND VGND VPWR VPWR _10512_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21020_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[27\] _02468_ VGND
+ VGND VPWR VPWR _02786_ sky130_fd_sc_hd__nand2_2
XFILLER_0_168_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22971_ _10583_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__buf_2
XFILLER_0_184_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_241_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21922_ _03453_ _03638_ _03619_ _03612_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_184_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_804 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24641_ clknet_leaf_22_clk net261 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[117\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21853_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[25\] _03376_ VGND
+ VGND VPWR VPWR _03573_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20804_ _02549_ _02578_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24572_ clknet_leaf_140_clk _01105_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dfxtp_4
X_21784_ _03484_ _03487_ _03506_ _01984_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23523_ clknet_leaf_138_clk _00056_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20735_ _02493_ _02511_ _07595_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23454_ net740 _04840_ _04849_ _04844_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20666_ _02444_ _02445_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22405_ _04005_ _04007_ _04046_ _04052_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__a31o_1
XFILLER_0_144_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23385_ net810 _04804_ _04812_ _04808_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__o211a_1
X_20597_ _02314_ _02340_ _02338_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_162_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22336_ _04020_ _04021_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22267_ _03953_ _03954_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_44_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24006_ clknet_leaf_46_clk _00539_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[7\]
+ sky130_fd_sc_hd__dfxtp_2
X_12020_ net816 _05018_ _05026_ _05022_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__o211a_1
XFILLER_0_218_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21218_ _02936_ _02939_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__nand2_1
X_22198_ _03880_ _03881_ _03886_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__a21o_2
XFILLER_0_44_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21149_ _02895_ _02021_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13971_ _06685_ _06689_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__xnor2_1
X_15710_ top_inst.grid_inst.data_path_wires\[7\]\[7\] _08149_ _08157_ _08154_ VGND
+ VGND VPWR VPWR _08326_ sky130_fd_sc_hd__nand4_1
X_12922_ _05658_ _05725_ _05656_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__o21ai_1
X_16690_ _09234_ _09235_ VGND VGND VPWR VPWR _09252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_214_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15641_ _08223_ _08224_ _08258_ VGND VGND VPWR VPWR _08259_ sky130_fd_sc_hd__a21o_1
XFILLER_0_213_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12853_ _05637_ _05619_ _05659_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__o21ai_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11804_ _04876_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__buf_2
XFILLER_0_51_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _10822_ _10824_ VGND VGND VPWR VPWR _10826_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15572_ _08191_ _08192_ VGND VGND VPWR VPWR _08193_ sky130_fd_sc_hd__and2_1
X_12784_ _05556_ _05558_ _05591_ _05592_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__a211oi_2
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[21\] _09628_ _09629_
+ VGND VGND VPWR VPWR _09854_ sky130_fd_sc_hd__a21oi_2
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14523_ _07213_ _07214_ net209 _07169_ VGND VGND VPWR VPWR _07216_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_16_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11735_ net35 net166 VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_132_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18291_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[7\] _10757_ VGND
+ VGND VPWR VPWR _10758_ sky130_fd_sc_hd__xor2_1
XFILLER_0_113_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_189_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17242_ _09761_ _09781_ VGND VGND VPWR VPWR _09788_ sky130_fd_sc_hd__nand2_1
X_14454_ _07146_ _07147_ _07145_ VGND VGND VPWR VPWR _07149_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_83_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13405_ _06170_ _06171_ _06176_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__o21a_1
X_17173_ _09707_ _09709_ VGND VGND VPWR VPWR _09722_ sky130_fd_sc_hd__and2_1
X_14385_ _07085_ VGND VGND VPWR VPWR _07086_ sky130_fd_sc_hd__buf_2
XFILLER_0_98_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16124_ _08667_ _08686_ _08664_ _08683_ VGND VGND VPWR VPWR _08712_ sky130_fd_sc_hd__nand4_1
X_13336_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[12\] _05354_ _06109_
+ _06110_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_5__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_4_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16055_ top_inst.grid_inst.data_path_wires\[8\]\[0\] VGND VGND VPWR VPWR _08661_
+ sky130_fd_sc_hd__buf_2
XFILLER_0_121_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13267_ top_inst.grid_inst.data_path_wires\[1\]\[4\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__and2b_1
XFILLER_0_84_1098 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15006_ _07649_ _07650_ VGND VGND VPWR VPWR _07660_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12218_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[2\] _05129_
+ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13198_ _05974_ _05975_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__xor2_1
XFILLER_0_62_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19814_ _01637_ _01639_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12149_ net398 _05097_ _05099_ _05088_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_236_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19745_ _01534_ _01571_ _01572_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__nand3_1
XFILLER_0_208_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16957_ _09360_ _09201_ net216 top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _09512_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_237_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15908_ _08149_ _08169_ _08518_ VGND VGND VPWR VPWR _08519_ sky130_fd_sc_hd__and3_1
X_19676_ _01476_ _01504_ _01505_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16888_ _09443_ _09444_ VGND VGND VPWR VPWR _09445_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_1014 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18627_ _11049_ _11050_ _11060_ _11058_ VGND VGND VPWR VPWR _11086_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15839_ _08374_ VGND VGND VPWR VPWR _08452_ sky130_fd_sc_hd__buf_4
XFILLER_0_232_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18558_ _10977_ _10979_ _11017_ VGND VGND VPWR VPWR _11019_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17509_ _10035_ _10033_ _10036_ _10024_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18489_ _10949_ _10951_ VGND VGND VPWR VPWR _10952_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_13 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20520_ _02301_ _02302_ _02271_ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_24 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_35 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_46 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_57 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20451_ _02226_ _02235_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__xnor2_1
XANTENNA_68 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_79 net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23170_ net799 _04685_ _04689_ _04691_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__o211a_1
X_20382_ _02129_ _02127_ _02125_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_207_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22121_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[5\] _03788_ _03789_
+ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput120 net120 VGND VGND VPWR VPWR output_tdata[59] sky130_fd_sc_hd__buf_2
XFILLER_0_140_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput131 net131 VGND VGND VPWR VPWR output_tdata[69] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput142 net142 VGND VGND VPWR VPWR output_tdata[79] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22052_ _03743_ _03744_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[3\]
+ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__a21oi_1
XTAP_6519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput153 net153 VGND VGND VPWR VPWR output_tdata[89] sky130_fd_sc_hd__buf_2
Xoutput164 net164 VGND VGND VPWR VPWR output_tdata[99] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21003_ _02768_ _02767_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__or2b_1
XTAP_5818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_242_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22954_ net389 _04557_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21905_ _03620_ _03621_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22885_ net708 _04522_ _04526_ _04524_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24624_ clknet_leaf_25_clk net372 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[100\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21836_ _03279_ _03556_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24555_ clknet_leaf_133_clk _01088_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21767_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[20\] _03421_ _03422_
+ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_194_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_1110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23506_ clknet_leaf_134_clk net455 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20718_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[15\] _02470_ VGND
+ VGND VPWR VPWR _02496_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24486_ clknet_leaf_84_clk net285 VGND VGND VPWR VPWR top_inst.valid_pipe\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21698_ _03279_ _03424_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23437_ _05736_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20649_ _02001_ _02227_ _02405_ _02406_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_191_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14170_ _06839_ _06841_ VGND VGND VPWR VPWR _06884_ sky130_fd_sc_hd__nor2_1
X_23368_ net833 _04791_ _04802_ _04795_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13121_ _05888_ _05900_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__xnor2_1
X_22319_ _03932_ _03930_ _03971_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23299_ net804 _04752_ _04763_ _04756_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__o211a_1
X_13052_ _05832_ _05833_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__nor2_1
XFILLER_0_237_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12003_ net894 _05004_ _05016_ _05008_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17860_ _10328_ _10331_ _10365_ VGND VGND VPWR VPWR _10366_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_100_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16811_ _09362_ _09368_ VGND VGND VPWR VPWR _09369_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_218_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17791_ top_inst.grid_inst.data_path_wires\[11\]\[2\] _10059_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[6\]
+ top_inst.grid_inst.data_path_wires\[11\]\[3\] VGND VGND VPWR VPWR _10299_ sky130_fd_sc_hd__and4b_1
XFILLER_0_206_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_13__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_4_13__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19530_ _11701_ _11692_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16742_ _09295_ _09300_ _09301_ VGND VGND VPWR VPWR _09302_ sky130_fd_sc_hd__nand3_2
X_13954_ _06624_ _06640_ _06637_ _06626_ VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12905_ _05682_ _05683_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__or2b_1
XFILLER_0_202_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16673_ _09233_ _09234_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[2\]
+ VGND VGND VPWR VPWR _09236_ sky130_fd_sc_hd__a21o_1
X_19461_ _11722_ _01295_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__and2_1
XFILLER_0_186_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13885_ _06622_ _06620_ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18412_ _10836_ _10876_ VGND VGND VPWR VPWR _10877_ sky130_fd_sc_hd__xnor2_1
X_12836_ _05639_ _05642_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_1032 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15624_ _08143_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[2\] _08240_
+ _08241_ VGND VGND VPWR VPWR _08242_ sky130_fd_sc_hd__a22o_1
X_19392_ _01197_ _01223_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__nor2_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15555_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[1\] _08175_ _08176_
+ VGND VGND VPWR VPWR _08177_ sky130_fd_sc_hd__nand3_1
X_18343_ _10806_ _10808_ VGND VGND VPWR VPWR _10809_ sky130_fd_sc_hd__xnor2_1
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _05574_ _05575_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _07196_ _07197_ _07191_ VGND VGND VPWR VPWR _07199_ sky130_fd_sc_hd__a21o_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18274_ _10739_ _10740_ _10711_ _10712_ VGND VGND VPWR VPWR _10742_ sky130_fd_sc_hd__o211ai_1
X_15486_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[15\] _07924_ _07844_
+ VGND VGND VPWR VPWR _08126_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12698_ _05506_ _05507_ _05508_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__or3_4
XFILLER_0_167_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17225_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[18\] _09631_ VGND
+ VGND VPWR VPWR _09772_ sky130_fd_sc_hd__xnor2_2
X_14437_ _07113_ _07132_ VGND VGND VPWR VPWR _07133_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput11 input_tdata[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_4
XFILLER_0_86_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput22 input_tdata[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput33 input_tvalid VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_4
XFILLER_0_25_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17156_ _09703_ _09705_ VGND VGND VPWR VPWR _09706_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14368_ top_inst.skew_buff_inst.row\[1\].output_reg\[3\] top_inst.axis_in_inst.inbuf_bus\[11\]
+ _05266_ VGND VGND VPWR VPWR _07072_ sky130_fd_sc_hd__mux2_4
Xhold806 top_inst.axis_out_inst.out_buff_data\[0\] VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ _08677_ _08681_ _08698_ _08692_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__o211a_1
Xhold817 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[10\] VGND
+ VGND VPWR VPWR net999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[10\] VGND VGND
+ VPWR VPWR net1010 sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ _06081_ _06056_ _06092_ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__nand3_1
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17087_ _09636_ _09637_ _09597_ VGND VGND VPWR VPWR _09639_ sky130_fd_sc_hd__a21o_1
Xhold839 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[12\] VGND
+ VGND VPWR VPWR net1021 sky130_fd_sc_hd__dlygate4sd3_1
X_14299_ _06936_ _06972_ _07008_ VGND VGND VPWR VPWR _07009_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_126_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16038_ _08642_ _08644_ VGND VGND VPWR VPWR _08646_ sky130_fd_sc_hd__nor2_1
XFILLER_0_204_1358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17989_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[14\] _10367_ VGND
+ VGND VPWR VPWR _10492_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_237_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19728_ _01518_ _01556_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__xor2_2
XFILLER_0_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19659_ _11701_ _11704_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__and2_1
XFILLER_0_215_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22670_ _04310_ _04343_ _04309_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21621_ _03210_ _03329_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24340_ clknet_leaf_8_clk _00873_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[99\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21552_ _03281_ _03283_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20503_ top_inst.grid_inst.data_path_wires\[16\]\[6\] top_inst.grid_inst.data_path_wires\[16\]\[5\]
+ _02013_ _02011_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__and4_1
X_24271_ clknet_leaf_97_clk _00804_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21483_ _02873_ _02893_ _03175_ _03216_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23222_ net513 _04713_ _04720_ _04717_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__o211a_1
X_20434_ net745 _01735_ _02219_ _02035_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_244_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23153_ net73 _04672_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__or2_1
X_20365_ _02149_ _02150_ _02151_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__nand3_1
XFILLER_0_113_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22104_ _03741_ _03761_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23084_ top_inst.axis_in_inst.inbuf_bus\[29\] _04629_ VGND VGND VPWR VPWR _04640_
+ sky130_fd_sc_hd__or2_1
X_20296_ _02083_ _02084_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__and2b_1
XTAP_6316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22035_ _03719_ _03720_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__nand2_1
XTAP_6349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23986_ clknet_leaf_80_clk _00519_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_242_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22937_ net621 _04543_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13670_ _06367_ _06370_ _06368_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__o21ba_1
X_22868_ net715 _04509_ _04516_ _04511_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12621_ _05432_ _05433_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__xor2_1
XFILLER_0_196_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24607_ clknet_leaf_25_clk _01140_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_116_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21819_ _03539_ _03540_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22799_ _04268_ _04431_ _04448_ _04452_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__o31a_1
XFILLER_0_38_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15340_ _07949_ _07984_ VGND VGND VPWR VPWR _07985_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_241_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12552_ _05284_ _05283_ _05363_ _05366_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__o2bb2a_1
X_24538_ clknet_leaf_101_clk _01071_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dfxtp_4
XPHY_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15271_ _07621_ _07635_ _07633_ top_inst.grid_inst.data_path_wires\[6\]\[7\] VGND
+ VGND VPWR VPWR _07917_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24469_ clknet_leaf_40_clk _01002_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_12483_ _05290_ _05301_ _05303_ _05261_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17010_ _09509_ net226 _09516_ VGND VGND VPWR VPWR _09564_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_136_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14222_ _06860_ _06898_ _06933_ VGND VGND VPWR VPWR _06934_ sky130_fd_sc_hd__nor3_1
XFILLER_0_22_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14153_ _06630_ _06648_ _06628_ _06645_ VGND VGND VPWR VPWR _06867_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_100_clk clknet_4_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_120_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13104_ _05352_ _05884_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__and2_1
X_14084_ _06738_ _06799_ _06758_ VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__a21oi_2
X_18961_ _11375_ _11377_ _11373_ VGND VGND VPWR VPWR _11383_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_954 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13035_ _05800_ _05817_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__nand2_1
X_17912_ _10415_ _10416_ VGND VGND VPWR VPWR _10417_ sky130_fd_sc_hd__nor2_1
X_18892_ top_inst.grid_inst.data_path_wires\[13\]\[0\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _11316_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17843_ _10332_ _10349_ VGND VGND VPWR VPWR _10350_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_206_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17774_ _10280_ _10281_ VGND VGND VPWR VPWR _10282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_221_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14986_ _07622_ _07639_ _07642_ _07643_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__o211a_1
XFILLER_0_234_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19513_ _01328_ _01330_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__nor2_1
X_16725_ _09253_ _09284_ _09285_ VGND VGND VPWR VPWR _09286_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_152_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13937_ net1000 _05403_ VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19444_ _01242_ _01277_ _01278_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__nand3_1
XFILLER_0_134_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16656_ _09189_ _09187_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _09221_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13868_ _06608_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12819_ _05547_ _05589_ _05587_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_201_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15607_ _08139_ _08159_ VGND VGND VPWR VPWR _08226_ sky130_fd_sc_hd__nand2_1
X_19375_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[2\] _11687_ VGND
+ VGND VPWR VPWR _01212_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16587_ _09135_ _09136_ _09133_ VGND VGND VPWR VPWR _09162_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13799_ _06541_ VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18326_ top_inst.grid_inst.data_path_wires\[12\]\[7\] _10600_ _10597_ VGND VGND VPWR
+ VPWR _10792_ sky130_fd_sc_hd__and3_1
XFILLER_0_151_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15538_ _08164_ _07641_ VGND VGND VPWR VPWR _08165_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15469_ _08101_ _08109_ VGND VGND VPWR VPWR _08110_ sky130_fd_sc_hd__xnor2_1
X_18257_ _10577_ _10612_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[5\]
+ _10599_ VGND VGND VPWR VPWR _10725_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_114_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17208_ _09753_ _09754_ _09623_ VGND VGND VPWR VPWR _09756_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_25_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18188_ _10642_ _10657_ _10658_ VGND VGND VPWR VPWR _10659_ sky130_fd_sc_hd__or3_1
Xhold603 _00930_ VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_887 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17139_ _09665_ _09689_ VGND VGND VPWR VPWR _09690_ sky130_fd_sc_hd__xor2_1
XFILLER_0_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold614 top_inst.axis_out_inst.out_buff_data\[50\] VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold625 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[10\] VGND
+ VGND VPWR VPWR net807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold636 top_inst.deskew_buff_inst.col_input\[77\] VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold647 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[11\] VGND
+ VGND VPWR VPWR net829 sky130_fd_sc_hd__dlygate4sd3_1
X_20150_ _01959_ _01960_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__or2_1
Xhold658 _00051_ VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold669 _00909_ VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20081_ _01893_ _01894_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23840_ clknet_leaf_89_clk _00373_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23771_ clknet_leaf_62_clk _00304_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20983_ _02749_ _02750_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__and2_1
XFILLER_0_240_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22722_ _04392_ _04393_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22653_ _04293_ _04327_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21604_ _03314_ _03334_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22584_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[18\] _04215_ _04216_
+ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__a21o_1
XFILLER_0_164_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24323_ clknet_leaf_5_clk _00856_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[18\]\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_111_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21535_ _03243_ _03267_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_895 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24254_ clknet_leaf_110_clk _00787_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21466_ _03163_ _03166_ _03199_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__a21bo_1
X_23205_ net676 _04700_ _04710_ _04704_ VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20417_ _02199_ _02200_ _02201_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__a21oi_1
X_24185_ clknet_leaf_47_clk _00718_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_21397_ _03132_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23136_ net165 _04659_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__or2_1
X_20348_ _04873_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__clkbuf_4
XTAP_6102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23067_ net1109 _04629_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__or2_1
XTAP_6146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20279_ _02066_ _02067_ _02050_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22018_ _03698_ _03680_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__and3_1
XTAP_6179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ _07523_ _07524_ VGND VGND VPWR VPWR _07525_ sky130_fd_sc_hd__nor2_1
XTAP_5478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14771_ _07417_ _07419_ VGND VGND VPWR VPWR _07458_ sky130_fd_sc_hd__nand2_1
XFILLER_0_192_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23969_ clknet_leaf_85_clk _00502_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_11983_ top_inst.axis_out_inst.out_buff_data\[61\] _04996_ VGND VGND VPWR VPWR _05005_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_242_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16510_ _09085_ _09086_ VGND VGND VPWR VPWR _09087_ sky130_fd_sc_hd__xnor2_1
X_13722_ _06385_ _06466_ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17490_ _05736_ _09187_ VGND VGND VPWR VPWR _10023_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16441_ _09018_ _09019_ VGND VGND VPWR VPWR _09020_ sky130_fd_sc_hd__or2b_1
XFILLER_0_128_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13653_ _06353_ _06354_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__or2b_1
XFILLER_0_195_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12604_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[3\]
+ _05282_ _05287_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__and4_1
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16372_ _08949_ _08951_ VGND VGND VPWR VPWR _08953_ sky130_fd_sc_hd__and2_1
X_19160_ _11576_ _11577_ VGND VGND VPWR VPWR _11578_ sky130_fd_sc_hd__or2_1
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13584_ _06330_ _06331_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15323_ _07952_ _07953_ _07967_ VGND VGND VPWR VPWR _07968_ sky130_fd_sc_hd__a21oi_1
X_18111_ _10038_ _10584_ _10593_ _10594_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12535_ _05349_ _05350_ _05336_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_152_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19091_ _11488_ _11490_ VGND VGND VPWR VPWR _11510_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15254_ _07898_ _07900_ VGND VGND VPWR VPWR _07901_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18042_ _10521_ _10519_ VGND VGND VPWR VPWR _10543_ sky130_fd_sc_hd__nand2_1
X_12466_ _05270_ _05287_ _05289_ _05261_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14205_ _06914_ _06916_ VGND VGND VPWR VPWR _06918_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15185_ _07619_ _07615_ _07635_ _07633_ VGND VGND VPWR VPWR _07833_ sky130_fd_sc_hd__nand4_4
XFILLER_0_201_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12397_ net323 _05235_ VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_238_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14136_ _06652_ _06626_ _06849_ VGND VGND VPWR VPWR _06850_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19993_ _01809_ _01810_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_238_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14067_ _06744_ _06746_ VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__nand2_1
X_18944_ _11322_ _11299_ VGND VGND VPWR VPWR _11367_ sky130_fd_sc_hd__or2b_1
XFILLER_0_201_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13018_ net1073 _05788_ _05801_ _05767_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18875_ _11271_ _11280_ _11282_ VGND VGND VPWR VPWR _11299_ sky130_fd_sc_hd__o21ai_1
XTAP_6680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17826_ _10304_ _10303_ VGND VGND VPWR VPWR _10333_ sky130_fd_sc_hd__or2b_1
XFILLER_0_206_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17757_ _10262_ _10265_ VGND VGND VPWR VPWR _10266_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_221_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14969_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _07631_ sky130_fd_sc_hd__buf_4
XFILLER_0_222_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16708_ _09207_ _09186_ net1120 _09203_ VGND VGND VPWR VPWR _09269_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17688_ _10037_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[0\]
+ top_inst.grid_inst.data_path_wires\[11\]\[7\] VGND VGND VPWR VPWR _10198_ sky130_fd_sc_hd__a22o_1
X_19427_ _11683_ net195 _11704_ _11678_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__a22o_1
X_16639_ _09207_ _09199_ VGND VGND VPWR VPWR _09208_ sky130_fd_sc_hd__or2_1
XFILLER_0_174_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19358_ _01182_ _01183_ _01194_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18309_ _10752_ _10775_ VGND VGND VPWR VPWR _10776_ sky130_fd_sc_hd__xor2_1
XFILLER_0_190_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19289_ _09185_ _11687_ _11690_ _11641_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21320_ _03043_ _03057_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold400 _01154_ VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__dlygate4sd3_1
X_21251_ _02135_ _02990_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__and2_1
XFILLER_0_241_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold411 _00178_ VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 top_inst.deskew_buff_inst.col_input\[68\] VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold433 _00022_ VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__dlygate4sd3_1
X_20202_ _02003_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__buf_4
Xhold444 _00007_ VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[6\] VGND VGND
+ VPWR VPWR net637 sky130_fd_sc_hd__dlygate4sd3_1
X_21182_ _02862_ _02889_ _02887_ _02864_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__a22o_1
XFILLER_0_180_1280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold466 top_inst.deskew_buff_inst.col_input\[85\] VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap174 _02360_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_1351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold477 top_inst.deskew_buff_inst.col_input\[108\] VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20133_ _01915_ _01922_ _01940_ _01896_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__a22oi_4
Xhold488 top_inst.deskew_buff_inst.col_input\[87\] VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[4\] VGND VGND
+ VPWR VPWR net681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20064_ _01853_ _01869_ _01878_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23823_ clknet_leaf_94_clk _00356_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23754_ clknet_leaf_135_clk net287 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1068 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20966_ _02733_ _02734_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__nand2_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22705_ _04365_ _04376_ _04367_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__or3_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23685_ clknet_leaf_118_clk _00218_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20897_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[21\] _02666_ _02667_
+ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__o21a_1
XFILLER_0_222_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22636_ _04307_ _04311_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__xor2_2
XFILLER_0_14_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22567_ _04245_ _04237_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__xor2_2
XFILLER_0_106_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24306_ clknet_leaf_138_clk _00839_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[81\]
+ sky130_fd_sc_hd__dfxtp_1
X_12320_ net567 _05196_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21518_ _03249_ _03250_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22498_ _04149_ _04179_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_224_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12251_ net437 _05151_ _05158_ _05155_ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__o211a_1
X_24237_ clknet_leaf_113_clk _00770_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21449_ _03167_ _03183_ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_181_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24168_ clknet_leaf_8_clk _00701_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_31_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12182_ net341 _05110_ _05118_ _05114_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23119_ net77 _04659_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__or2_1
XFILLER_0_236_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16990_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[10\] _09459_ _09417_
+ VGND VGND VPWR VPWR _09544_ sky130_fd_sc_hd__a21o_1
X_24099_ clknet_leaf_15_clk _00632_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15941_ _08549_ _08551_ VGND VGND VPWR VPWR _08552_ sky130_fd_sc_hd__nor2_1
XFILLER_0_235_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18660_ _11109_ _11111_ VGND VGND VPWR VPWR _11117_ sky130_fd_sc_hd__nor2_1
XFILLER_0_244_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ _08409_ _08483_ VGND VGND VPWR VPWR _08484_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_235_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17611_ _10121_ _10122_ _09292_ VGND VGND VPWR VPWR _10124_ sky130_fd_sc_hd__a21o_1
X_14823_ _07467_ _07470_ _07508_ VGND VGND VPWR VPWR _07509_ sky130_fd_sc_hd__a21o_1
XFILLER_0_162_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18591_ _11049_ _11050_ VGND VGND VPWR VPWR _11051_ sky130_fd_sc_hd__nand2_1
XFILLER_0_230_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ _10059_ _10057_ VGND VGND VPWR VPWR _10060_ sky130_fd_sc_hd__or2_1
X_14754_ _07437_ _07359_ VGND VGND VPWR VPWR _07441_ sky130_fd_sc_hd__and2b_1
X_11966_ net805 _04990_ _04993_ _04995_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__o211a_1
XFILLER_0_230_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13705_ top_inst.grid_inst.data_path_wires\[2\]\[3\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__and2b_1
X_14685_ _07079_ _07086_ _07090_ _07074_ VGND VGND VPWR VPWR _07374_ sky130_fd_sc_hd__a22o_1
X_17473_ _09998_ _10007_ VGND VGND VPWR VPWR _10009_ sky130_fd_sc_hd__or2_1
X_11897_ _04876_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_1118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19212_ _11387_ _11590_ _11626_ VGND VGND VPWR VPWR _11628_ sky130_fd_sc_hd__nor3_1
XFILLER_0_156_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16424_ _08965_ _08964_ VGND VGND VPWR VPWR _09003_ sky130_fd_sc_hd__or2b_1
X_13636_ _06380_ _06382_ VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_776 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19143_ _11559_ _11560_ VGND VGND VPWR VPWR _11561_ sky130_fd_sc_hd__and2_1
XFILLER_0_172_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16355_ _08883_ _08886_ _08887_ _08935_ _08880_ VGND VGND VPWR VPWR _08936_ sky130_fd_sc_hd__a32oi_4
X_13567_ _06290_ _06291_ _06314_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__and3_1
XFILLER_0_165_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12518_ _05311_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__buf_8
X_15306_ _07933_ _07934_ VGND VGND VPWR VPWR _07951_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19074_ _11492_ _11493_ VGND VGND VPWR VPWR _11494_ sky130_fd_sc_hd__xnor2_1
X_16286_ _08831_ _08868_ VGND VGND VPWR VPWR _08869_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13498_ _06247_ _06248_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_1242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18025_ _10525_ _10526_ VGND VGND VPWR VPWR _10527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12449_ _05275_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__buf_4
X_15237_ _07830_ VGND VGND VPWR VPWR _07884_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15168_ _07814_ _07815_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[7\]
+ _07816_ VGND VGND VPWR VPWR _07817_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_10_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14119_ _06769_ _06781_ VGND VGND VPWR VPWR _06834_ sky130_fd_sc_hd__nand2_1
XFILLER_0_239_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19976_ _01754_ _01793_ _01794_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__a21o_1
X_15099_ top_inst.grid_inst.data_path_wires\[6\]\[3\] _07610_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _07749_ sky130_fd_sc_hd__nand4_4
XFILLER_0_61_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18927_ top_inst.grid_inst.data_path_wires\[13\]\[1\] top_inst.grid_inst.data_path_wires\[13\]\[2\]
+ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _11350_ sky130_fd_sc_hd__and4b_1
XFILLER_0_24_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18858_ _11270_ _11281_ VGND VGND VPWR VPWR _11283_ sky130_fd_sc_hd__or2_1
X_17809_ _10314_ _10316_ VGND VGND VPWR VPWR _10317_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18789_ _11214_ _11215_ VGND VGND VPWR VPWR _11216_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20820_ _02593_ _02590_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20751_ _02517_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23470_ clknet_leaf_32_clk net565 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[124\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20682_ _02364_ _02440_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__and2_1
XFILLER_0_174_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22421_ _03711_ _03693_ _04068_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__and3_1
XFILLER_0_169_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_843 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22352_ _04022_ _04037_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__xor2_2
XFILLER_0_198_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21303_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[7\] _03040_ VGND
+ VGND VPWR VPWR _03041_ sky130_fd_sc_hd__xor2_2
XFILLER_0_108_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_1315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22283_ _03969_ _03970_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_1435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24022_ clknet_leaf_55_clk _00555_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold230 _00055_ VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__dlygate4sd3_1
X_21234_ top_inst.grid_inst.data_path_wires\[17\]\[4\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[1\]
+ _02882_ top_inst.grid_inst.data_path_wires\[17\]\[5\] VGND VGND VPWR VPWR _02974_
+ sky130_fd_sc_hd__a22o_1
Xhold241 top_inst.axis_out_inst.out_buff_data\[110\] VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold252 top_inst.axis_out_inst.out_buff_data\[92\] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[8\] VGND
+ VGND VPWR VPWR net445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[3\] VGND
+ VGND VPWR VPWR net456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold285 top_inst.axis_out_inst.out_buff_enabled VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21165_ _02706_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_217_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold296 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[3\] VGND
+ VGND VPWR VPWR net478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1083 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20116_ _01927_ _01928_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21096_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[27\] _02666_ VGND
+ VGND VPWR VPWR _02858_ sky130_fd_sc_hd__and2b_1
XFILLER_0_233_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_217_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20047_ _07707_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_232_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_1400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11820_ _04911_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__clkbuf_4
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _05275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23806_ clknet_leaf_76_clk _00339_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA_114 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21998_ _02706_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__clkbuf_4
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11751_ net630 _04860_ _04871_ _04870_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__o211a_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23737_ clknet_leaf_127_clk _00270_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_20949_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[24\] _02468_ VGND
+ VGND VPWR VPWR _02718_ sky130_fd_sc_hd__nand2_1
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_80_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14470_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[0\]
+ _07077_ _07081_ VGND VGND VPWR VPWR _07164_ sky130_fd_sc_hd__nand4_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23668_ clknet_leaf_125_clk net409 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13421_ _06188_ _05262_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22619_ _04271_ _04286_ _04295_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23599_ clknet_leaf_103_clk net328 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16140_ _08724_ _08726_ VGND VGND VPWR VPWR _08727_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13352_ _06090_ _06089_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__or2b_1
XFILLER_0_84_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12303_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[6\] _05183_
+ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16071_ _08163_ _08663_ _08672_ _08666_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__o211a_1
X_13283_ _06014_ _06013_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__and2b_1
XFILLER_0_161_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15022_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[3\] _07673_ _07674_
+ VGND VGND VPWR VPWR _07675_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12234_ net846 _05137_ _05148_ _05141_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19830_ _01562_ _01634_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12165_ net592 _05097_ _05108_ _05101_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19761_ _01522_ _01549_ _01548_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_159_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16973_ _09525_ _09526_ _09499_ VGND VGND VPWR VPWR _09528_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12096_ net272 _05058_ _05069_ _05062_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18712_ _11149_ _11150_ VGND VGND VPWR VPWR _11151_ sky130_fd_sc_hd__or2_1
XTAP_5050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15924_ _08532_ _08533_ VGND VGND VPWR VPWR _08535_ sky130_fd_sc_hd__and2_1
XTAP_5061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19692_ _01481_ _01479_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__and2b_1
XFILLER_0_235_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 input_tdata[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XTAP_5083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18643_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[15\] _10923_ _10840_
+ VGND VGND VPWR VPWR _11101_ sky130_fd_sc_hd__a21o_1
XTAP_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _08429_ _08466_ VGND VGND VPWR VPWR _08468_ sky130_fd_sc_hd__nor2_1
XTAP_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ _07487_ _07491_ VGND VGND VPWR VPWR _07492_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18574_ _11033_ _11034_ VGND VGND VPWR VPWR _11035_ sky130_fd_sc_hd__and2_1
XFILLER_0_235_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15786_ _08398_ _08399_ VGND VGND VPWR VPWR _08400_ sky130_fd_sc_hd__nor2_1
XFILLER_0_231_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12998_ _05781_ _05782_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17525_ _10047_ _09199_ VGND VGND VPWR VPWR _10048_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14737_ _07410_ _07411_ _07424_ VGND VGND VPWR VPWR _07425_ sky130_fd_sc_hd__a21o_1
XFILLER_0_197_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11949_ net913 _04977_ _04985_ _04981_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_71_clk clknet_4_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_143_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17456_ _09980_ _09982_ VGND VGND VPWR VPWR _09992_ sky130_fd_sc_hd__or2b_1
XFILLER_0_15_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14668_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[9\] _07048_ _07356_
+ _07357_ _06180_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__o221a_1
XFILLER_0_172_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16407_ _08944_ _08946_ VGND VGND VPWR VPWR _08987_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13619_ top_inst.grid_inst.data_path_wires\[2\]\[1\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17387_ _09908_ _09909_ _09926_ VGND VGND VPWR VPWR _09927_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14599_ _07068_ VGND VGND VPWR VPWR _07290_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19126_ _11505_ _11543_ VGND VGND VPWR VPWR _11545_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16338_ _08872_ _08916_ _08914_ VGND VGND VPWR VPWR _08919_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_242_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19057_ _11158_ _11156_ _11147_ VGND VGND VPWR VPWR _11477_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_42_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16269_ _08849_ _08850_ _08801_ _08803_ VGND VGND VPWR VPWR _08852_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18008_ _10488_ _10510_ VGND VGND VPWR VPWR _10511_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19959_ _01763_ _01768_ _01766_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__a21o_1
XFILLER_0_215_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22970_ net718 _04562_ _04574_ _04564_ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__o211a_1
XFILLER_0_241_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21921_ _03598_ _03617_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__nand2_1
XFILLER_0_218_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24640_ clknet_leaf_25_clk net534 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[116\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21852_ _03555_ _03558_ _03557_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_195_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20803_ _02576_ _02577_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24571_ clknet_leaf_143_clk _01104_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21783_ _03484_ _03487_ _03506_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_62_clk clknet_4_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_16
X_23522_ clknet_leaf_139_clk net412 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1062 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20734_ _02493_ _02511_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23453_ net725 _04864_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20665_ _02426_ _02427_ _02443_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__and3_1
XFILLER_0_162_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22404_ _03070_ _04087_ _04088_ _03929_ VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23384_ net55 _04805_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__or2_1
X_20596_ _02354_ _02377_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_225_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22335_ _04016_ _04019_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22266_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[18\]\[3\]
+ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24005_ clknet_leaf_46_clk _00538_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_44_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21217_ _02955_ _02957_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__xor2_2
XFILLER_0_143_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22197_ _03838_ _03879_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__nor2_1
XFILLER_0_218_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21148_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _02895_ sky130_fd_sc_hd__buf_2
XFILLER_0_218_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13970_ _06670_ _06688_ VGND VGND VPWR VPWR _06689_ sky130_fd_sc_hd__xor2_1
X_21079_ _02643_ _02841_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_1040 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12921_ _05708_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__inv_2
XFILLER_0_244_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15640_ _08201_ _08222_ VGND VGND VPWR VPWR _08258_ sky130_fd_sc_hd__nor2_1
XFILLER_0_244_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12852_ _05653_ _05658_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11803_ net614 _04898_ _04901_ _04902_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__o211a_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _05562_ _05554_ _05590_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__and3_1
X_15571_ _08189_ _08190_ VGND VGND VPWR VPWR _08192_ sky130_fd_sc_hd__nand2_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_53_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_150_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _09834_ _09837_ _09836_ VGND VGND VPWR VPWR _09853_ sky130_fd_sc_hd__a21bo_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ net209 _07169_ _07213_ _07214_ VGND VGND VPWR VPWR _07215_ sky130_fd_sc_hd__a211o_1
XFILLER_0_138_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11734_ top_inst.axis_in_inst.inbuf_valid _04856_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__nand2_8
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18290_ _10755_ _10756_ VGND VGND VPWR VPWR _10757_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17241_ _05406_ VGND VGND VPWR VPWR _09787_ sky130_fd_sc_hd__buf_6
XFILLER_0_83_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14453_ _07145_ _07146_ _07147_ VGND VGND VPWR VPWR _07148_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_148_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13404_ _06172_ _06175_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14384_ top_inst.skew_buff_inst.row\[1\].output_reg\[6\] top_inst.axis_in_inst.inbuf_bus\[14\]
+ net208 VGND VGND VPWR VPWR _07085_ sky130_fd_sc_hd__mux2_4
X_17172_ _09583_ _09662_ _09718_ _09719_ _09720_ VGND VGND VPWR VPWR _09721_ sky130_fd_sc_hd__o311a_4
XFILLER_0_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13335_ _06080_ _06077_ _06108_ _05405_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__a31oi_1
X_16123_ _08686_ _08664_ _08683_ _08667_ VGND VGND VPWR VPWR _08711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13266_ _06035_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__inv_2
X_16054_ _06848_ _08659_ _08660_ _08166_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15005_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[2\] _07658_ VGND
+ VGND VPWR VPWR _07659_ sky130_fd_sc_hd__xor2_1
XFILLER_0_122_1218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12217_ net932 _05137_ _05138_ _05128_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13197_ _05927_ _05930_ _05928_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_161_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19813_ _01604_ _01632_ _01638_ _01613_ _01603_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__a32o_1
XFILLER_0_236_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12148_ top_inst.axis_out_inst.out_buff_data\[4\] _05089_ VGND VGND VPWR VPWR _05099_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_97_1416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19744_ _01298_ _11705_ _11708_ _11703_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__a2bb2o_1
X_16956_ _09360_ _09377_ _09201_ net227 VGND VGND VPWR VPWR _09511_ sky130_fd_sc_hd__or4b_4
X_12079_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[6\] _05050_
+ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__or2_1
XFILLER_0_223_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15907_ _08147_ _08353_ VGND VGND VPWR VPWR _08518_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19675_ _01502_ _01503_ _01456_ _01477_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_223_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16887_ _09441_ _09442_ _09386_ _09388_ VGND VGND VPWR VPWR _09444_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18626_ _11077_ _11084_ VGND VGND VPWR VPWR _11085_ sky130_fd_sc_hd__xor2_1
XFILLER_0_189_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15838_ _08449_ _08450_ VGND VGND VPWR VPWR _08451_ sky130_fd_sc_hd__nor2_1
XFILLER_0_220_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18557_ _10977_ _10979_ _11017_ VGND VGND VPWR VPWR _11018_ sky130_fd_sc_hd__o21ai_1
X_15769_ _08323_ _08332_ _08383_ VGND VGND VPWR VPWR _08384_ sky130_fd_sc_hd__o21a_1
XFILLER_0_188_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17508_ _10030_ _09210_ VGND VGND VPWR VPWR _10036_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18488_ _10907_ _10908_ _10950_ VGND VGND VPWR VPWR _10951_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17439_ _09974_ _09975_ VGND VGND VPWR VPWR _09976_ sky130_fd_sc_hd__nand2_1
XANTENNA_14 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_25 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_47 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20450_ _02228_ _02234_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__xnor2_1
XANTENNA_69 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19109_ _11526_ _11527_ VGND VGND VPWR VPWR _11528_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20381_ _02166_ _02167_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__or2_2
XFILLER_0_3_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22120_ _03785_ _03793_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput110 net110 VGND VGND VPWR VPWR output_tdata[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_203_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput121 net121 VGND VGND VPWR VPWR output_tdata[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput132 net132 VGND VGND VPWR VPWR output_tdata[6] sky130_fd_sc_hd__buf_2
Xoutput143 net143 VGND VGND VPWR VPWR output_tdata[7] sky130_fd_sc_hd__clkbuf_4
X_22051_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[3\] _03743_ _03744_
+ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__and3_1
XTAP_6509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput154 net154 VGND VGND VPWR VPWR output_tdata[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput165 net165 VGND VGND VPWR VPWR output_tdata[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21002_ _02767_ _02768_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__or2b_1
XFILLER_0_220_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22953_ net681 _04562_ _04565_ _04564_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21904_ _03620_ _03621_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__nor2_1
XFILLER_0_190_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22884_ top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[7\] _04517_ VGND
+ VGND VPWR VPWR _04526_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24623_ clknet_leaf_23_clk _01156_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[99\]
+ sky130_fd_sc_hd__dfxtp_1
X_21835_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[24\] _03376_ VGND
+ VGND VPWR VPWR _03556_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_clk clknet_4_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_210_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24554_ clknet_leaf_133_clk _01087_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_109_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21766_ _03473_ _03476_ _03475_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_182_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23505_ clknet_leaf_134_clk net429 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[95\]
+ sky130_fd_sc_hd__dfxtp_1
X_20717_ _02464_ _02475_ _02472_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__a21oi_1
X_24485_ clknet_leaf_115_clk _01018_ VGND VGND VPWR VPWR top_inst.valid_pipe\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21697_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[18\] _03376_ VGND
+ VGND VPWR VPWR _03424_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_230_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23436_ net893 _04827_ _04839_ _04831_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20648_ _02398_ _02400_ _02397_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23367_ net47 _04792_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20579_ _02359_ net174 VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_225_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13120_ _05894_ _05899_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22318_ _03969_ _04004_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__xor2_2
XFILLER_0_104_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23298_ net141 _04753_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__or2_1
XFILLER_0_221_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13051_ top_inst.grid_inst.data_path_wires\[1\]\[4\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[1\]\[5\]
+ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_131_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22249_ _03894_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12002_ net797 _05010_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__or2_1
XFILLER_0_218_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16810_ _09363_ _09367_ VGND VGND VPWR VPWR _09368_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_233_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17790_ _10032_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[5\] VGND
+ VGND VPWR VPWR _10298_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16741_ _09298_ _09299_ _09268_ _09270_ VGND VGND VPWR VPWR _09301_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_205_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13953_ _06661_ _06672_ VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__nand2_1
XFILLER_0_221_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12904_ _05658_ _05708_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__xor2_1
X_19460_ top_inst.deskew_buff_inst.col_input\[6\] _01294_ _08307_ VGND VGND VPWR VPWR
+ _01295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_236_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16672_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[2\] _09233_ _09234_
+ VGND VGND VPWR VPWR _09235_ sky130_fd_sc_hd__nand3_1
X_13884_ top_inst.grid_inst.data_path_wires\[3\]\[1\] VGND VGND VPWR VPWR _06622_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18411_ _10874_ _10875_ VGND VGND VPWR VPWR _10876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15623_ top_inst.grid_inst.data_path_wires\[7\]\[2\] top_inst.grid_inst.data_path_wires\[7\]\[1\]
+ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _08241_ sky130_fd_sc_hd__nand4_4
XFILLER_0_213_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12835_ _05447_ _05449_ _05297_ _05641_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__or4_1
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19391_ net812 _05634_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_clk clknet_4_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _10581_ _10610_ _10770_ _10807_ VGND VGND VPWR VPWR _10808_ sky130_fd_sc_hd__a31oi_2
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15554_ _08137_ _08135_ _08157_ _08155_ VGND VGND VPWR VPWR _08176_ sky130_fd_sc_hd__nand4_2
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12766_ _05293_ _05288_ _05301_ _05306_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__and4_1
XFILLER_0_185_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14505_ _07191_ _07196_ _07197_ VGND VGND VPWR VPWR _07198_ sky130_fd_sc_hd__nand3_2
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _10711_ _10712_ _10739_ _10740_ VGND VGND VPWR VPWR _10741_ sky130_fd_sc_hd__a211o_1
X_12697_ _05280_ _05273_ _05305_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__and3_1
X_15485_ _08107_ _08124_ VGND VGND VPWR VPWR _08125_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17224_ _09588_ _09753_ VGND VGND VPWR VPWR _09771_ sky130_fd_sc_hd__and2_1
X_14436_ _07130_ _07131_ VGND VGND VPWR VPWR _07132_ sky130_fd_sc_hd__and2b_1
Xinput12 input_tdata[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_114_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput23 input_tdata[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_8
Xinput34 load_weight VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_12
XFILLER_0_128_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17155_ _09623_ _09704_ VGND VGND VPWR VPWR _09705_ sky130_fd_sc_hd__xor2_1
X_14367_ _05290_ _07069_ _07071_ _06684_ VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold807 top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[31\] VGND VGND
+ VPWR VPWR net989 sky130_fd_sc_hd__dlygate4sd3_1
X_16106_ _08697_ _08684_ VGND VGND VPWR VPWR _08698_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold818 top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[1\] VGND VGND
+ VPWR VPWR net1000 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ _06081_ _06056_ _06092_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__a21o_1
XFILLER_0_204_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17086_ _09597_ _09636_ _09637_ VGND VGND VPWR VPWR _09638_ sky130_fd_sc_hd__nand3_1
X_14298_ _06971_ _06970_ VGND VGND VPWR VPWR _07008_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold829 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[13\] VGND VGND
+ VPWR VPWR net1011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16037_ _08620_ _08621_ _08618_ VGND VGND VPWR VPWR _08645_ sky130_fd_sc_hd__a21oi_1
X_13249_ _05945_ _06024_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17988_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[14\] _10367_ VGND
+ VGND VPWR VPWR _10491_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_1346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19727_ _01554_ _01555_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__nand2_2
X_16939_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[9\] _09494_ VGND
+ VGND VPWR VPWR _09495_ sky130_fd_sc_hd__or2_1
XFILLER_0_237_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19658_ _01486_ _01487_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__nand2_2
X_18609_ _11065_ _11068_ VGND VGND VPWR VPWR _11069_ sky130_fd_sc_hd__xor2_2
XFILLER_0_94_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19589_ _01418_ _01419_ net249 VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_clk clknet_4_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_1155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21620_ _03320_ _03331_ VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__and2b_1
XFILLER_0_133_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21551_ _03245_ _03282_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__xor2_1
XFILLER_0_168_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20502_ _02284_ _02285_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__xor2_2
XFILLER_0_133_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24270_ clknet_leaf_100_clk _00803_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_21482_ top_inst.grid_inst.data_path_wires\[17\]\[4\] _02895_ _03173_ VGND VGND VPWR
+ VPWR _03216_ sky130_fd_sc_hd__and3_1
XFILLER_0_173_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23221_ net104 _04714_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20433_ _05317_ _02218_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23152_ net955 _04671_ _04679_ _04675_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__o211a_1
X_20364_ top_inst.grid_inst.data_path_wires\[16\]\[4\] top_inst.grid_inst.data_path_wires\[16\]\[3\]
+ _02013_ _02051_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__nand4_2
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22103_ _03778_ _03794_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__xor2_2
XFILLER_0_12_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23083_ net21 _04628_ _04639_ _04632_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__o211a_1
XTAP_6306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20295_ _02081_ _02082_ _02077_ _02054_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22034_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[2\] _03728_ VGND
+ VGND VPWR VPWR _03729_ sky130_fd_sc_hd__xnor2_1
XTAP_6339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23985_ clknet_leaf_80_clk _00518_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_243_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22936_ net1007 _04548_ _04555_ _04551_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22867_ top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[0\] _04504_ VGND
+ VGND VPWR VPWR _04516_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12620_ _05384_ _05387_ _05388_ _05358_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__a22o_1
X_24606_ clknet_leaf_25_clk _01139_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_52_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21818_ _03537_ _03538_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__and2_1
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22798_ _04454_ _04455_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__or2b_1
XFILLER_0_116_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12551_ _05364_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24537_ clknet_leaf_129_clk _01070_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dfxtp_4
X_21749_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[20\] _03376_ VGND
+ VGND VPWR VPWR _03474_ sky130_fd_sc_hd__xnor2_1
XPHY_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_241_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12482_ _05302_ _05294_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__or2_1
XFILLER_0_191_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15270_ top_inst.grid_inst.data_path_wires\[6\]\[7\] _07635_ _07633_ VGND VGND VPWR
+ VPWR _07916_ sky130_fd_sc_hd__and3_1
X_24468_ clknet_leaf_54_clk _01001_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14221_ _06648_ _06645_ _06635_ VGND VGND VPWR VPWR _06933_ sky130_fd_sc_hd__o21ai_1
X_23419_ net1107 _04596_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__or2_1
X_24399_ clknet_leaf_38_clk _00932_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14152_ _06862_ _06865_ VGND VGND VPWR VPWR _06866_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13103_ _05881_ _05883_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[6\]
+ _05327_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__a2bb2o_1
X_14083_ _06756_ VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__inv_2
XFILLER_0_162_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18960_ _11366_ _11369_ VGND VGND VPWR VPWR _11382_ sky130_fd_sc_hd__nor2_1
XFILLER_0_237_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13034_ _05795_ _05816_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__xor2_1
X_17911_ _10412_ _10414_ VGND VGND VPWR VPWR _10416_ sky130_fd_sc_hd__and2_1
XFILLER_0_197_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18891_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[13\]\[1\]
+ VGND VGND VPWR VPWR _11315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17842_ _10347_ _10348_ VGND VGND VPWR VPWR _10349_ sky130_fd_sc_hd__or2_1
XFILLER_0_219_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1070 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17773_ _10232_ _10238_ VGND VGND VPWR VPWR _10281_ sky130_fd_sc_hd__or2b_1
XFILLER_0_206_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14985_ _07617_ VGND VGND VPWR VPWR _07643_ sky130_fd_sc_hd__clkbuf_4
X_19512_ _01339_ _01341_ _01338_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_135_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16724_ _09251_ _09252_ VGND VGND VPWR VPWR _09285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13936_ _05406_ _06656_ _06657_ VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__or3b_1
XFILLER_0_18_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19443_ _01272_ _01273_ _01276_ VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__a21o_1
X_16655_ net1058 _05276_ _09220_ _09184_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__o211a_1
X_13867_ _06364_ _06607_ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15606_ _08223_ _08224_ VGND VGND VPWR VPWR _08225_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_215_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12818_ _05624_ _05625_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19374_ _01207_ _01208_ _01209_ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16586_ _09159_ _09160_ VGND VGND VPWR VPWR _09161_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13798_ _06539_ _06540_ VGND VGND VPWR VPWR _06541_ sky130_fd_sc_hd__nand2_2
XFILLER_0_139_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18325_ _10600_ _10597_ top_inst.grid_inst.data_path_wires\[12\]\[7\] VGND VGND VPWR
+ VPWR _10791_ sky130_fd_sc_hd__o21ai_2
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15537_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _08164_ sky130_fd_sc_hd__clkbuf_4
X_12749_ _05556_ _05557_ _05520_ _05522_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__a211o_1
XFILLER_0_173_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18256_ _10684_ _10689_ VGND VGND VPWR VPWR _10724_ sky130_fd_sc_hd__or2b_1
XFILLER_0_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15468_ _08107_ _08108_ VGND VGND VPWR VPWR _08109_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17207_ _09623_ _09753_ _09754_ VGND VGND VPWR VPWR _09755_ sky130_fd_sc_hd__nand3b_1
X_14419_ _06364_ _07115_ VGND VGND VPWR VPWR _07116_ sky130_fd_sc_hd__and2_1
XFILLER_0_181_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18187_ _10643_ _10635_ _10655_ VGND VGND VPWR VPWR _10658_ sky130_fd_sc_hd__and3_1
X_15399_ _08030_ _07998_ _08040_ VGND VGND VPWR VPWR _08042_ sky130_fd_sc_hd__nand3_1
XFILLER_0_25_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17138_ _09666_ _09688_ VGND VGND VPWR VPWR _09689_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold604 top_inst.deskew_buff_inst.col_input\[24\] VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold615 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[5\] VGND
+ VGND VPWR VPWR net797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 top_inst.deskew_buff_inst.col_input\[72\] VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold637 _00052_ VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold648 top_inst.axis_out_inst.out_buff_data\[19\] VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__dlygate4sd3_1
X_17069_ _09583_ _09618_ _09616_ VGND VGND VPWR VPWR _09621_ sky130_fd_sc_hd__o21ai_1
Xhold659 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[10\] VGND
+ VGND VPWR VPWR net841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_6_clk clknet_4_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_16
X_20080_ _01562_ _01892_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__nand2_1
XFILLER_0_244_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23770_ clknet_leaf_62_clk _00303_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_20982_ _02528_ _02741_ _02748_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__nand3_1
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_1299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22721_ _04390_ _04391_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22652_ _04137_ _04312_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21603_ _03332_ _03333_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__xnor2_2
X_22583_ _04240_ _04243_ _04242_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21534_ _03265_ _03266_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__xnor2_1
X_24322_ clknet_leaf_10_clk _00855_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[18\]\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_209_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24253_ clknet_leaf_106_clk _00786_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21465_ _03165_ _03164_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__or2b_1
XFILLER_0_90_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23204_ net96 _04701_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20416_ _02199_ _02200_ _02201_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24184_ clknet_leaf_29_clk _00717_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21396_ top_inst.grid_inst.data_path_wires\[17\]\[6\] top_inst.grid_inst.data_path_wires\[17\]\[5\]
+ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__and4_1
X_23135_ net310 _04656_ _04669_ _04662_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__o211a_1
X_20347_ _05440_ _02134_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23066_ net13 _04628_ _04630_ _04619_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20278_ _02050_ _02066_ _02067_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__or3_4
XFILLER_0_235_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22017_ _03695_ _05270_ _03714_ _03702_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__o211a_1
XTAP_6169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_243_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14770_ _07415_ _07423_ VGND VGND VPWR VPWR _07457_ sky130_fd_sc_hd__nand2_1
XTAP_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ _04911_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__clkbuf_4
X_23968_ clknet_leaf_86_clk _00501_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_13721_ _06418_ _06421_ _06419_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__o21ba_1
X_22919_ net380 _04535_ _04545_ _04537_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23899_ clknet_leaf_52_clk _00432_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_808 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16440_ _09003_ _09004_ _09017_ VGND VGND VPWR VPWR _09019_ sky130_fd_sc_hd__nand3_1
XFILLER_0_79_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13652_ _06396_ _06398_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1085 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12603_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[4\] _05282_ _05287_
+ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _05416_ sky130_fd_sc_hd__a22oi_1
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16371_ _08949_ _08951_ VGND VGND VPWR VPWR _08952_ sky130_fd_sc_hd__nor2_1
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13583_ _06186_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[5\] VGND
+ VGND VPWR VPWR _06331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18110_ _10447_ VGND VGND VPWR VPWR _10594_ sky130_fd_sc_hd__clkbuf_4
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15322_ _07965_ _07966_ VGND VGND VPWR VPWR _07967_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12534_ _05347_ _05348_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__and2_1
X_19090_ _11508_ VGND VGND VPWR VPWR _11509_ sky130_fd_sc_hd__inv_2
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18041_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[15\] _08183_ _10542_
+ _10448_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__o211a_1
X_15253_ _07856_ _07857_ _07899_ VGND VGND VPWR VPWR _07900_ sky130_fd_sc_hd__o21a_1
X_12465_ _05288_ _05276_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14204_ _06914_ _06916_ VGND VGND VPWR VPWR _06917_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15184_ _07615_ _07635_ _07633_ _07619_ VGND VGND VPWR VPWR _07832_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12396_ net515 _05230_ _05240_ _05234_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14135_ top_inst.grid_inst.data_path_wires\[3\]\[2\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _06849_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19992_ _01800_ _01808_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_1170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14066_ _06769_ _06781_ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__xnor2_2
X_18943_ _11335_ _11365_ VGND VGND VPWR VPWR _11366_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_238_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13017_ _05799_ _05800_ _05336_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18874_ _11264_ _11268_ _11297_ VGND VGND VPWR VPWR _11298_ sky130_fd_sc_hd__o21ai_2
XTAP_6670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17825_ _10328_ _10331_ VGND VGND VPWR VPWR _10332_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17756_ _10263_ _10264_ VGND VGND VPWR VPWR _10265_ sky130_fd_sc_hd__and2_1
X_14968_ _07608_ _06647_ _07630_ _07618_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_234_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16707_ _09207_ _09203_ _09186_ net1120 VGND VGND VPWR VPWR _09268_ sky130_fd_sc_hd__nand4_4
XFILLER_0_7_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13919_ _06626_ _06204_ _06646_ _06639_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__o211a_1
X_17687_ _10172_ _10173_ VGND VGND VPWR VPWR _10197_ sky130_fd_sc_hd__nor2_1
X_14899_ _07531_ _07528_ VGND VGND VPWR VPWR _07582_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19426_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[5\] _01230_ _01231_
+ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_230_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16638_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _09207_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19357_ _01182_ _01183_ _01194_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__a21oi_2
X_16569_ _09143_ _09144_ VGND VGND VPWR VPWR _09145_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18308_ _10760_ _10774_ VGND VGND VPWR VPWR _10775_ sky130_fd_sc_hd__xnor2_1
X_19288_ _11688_ _11689_ VGND VGND VPWR VPWR _11690_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18239_ _10682_ _10706_ _08265_ VGND VGND VPWR VPWR _10708_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21250_ top_inst.deskew_buff_inst.col_input\[69\] _11723_ _02988_ _02989_ VGND VGND
+ VPWR VPWR _02990_ sky130_fd_sc_hd__a22o_1
Xhold401 top_inst.axis_in_inst.inbuf_bus\[14\] VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold412 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[3\] VGND
+ VGND VPWR VPWR net594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold423 top_inst.valid_pipe\[2\] VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__dlygate4sd3_1
X_20201_ top_inst.grid_inst.data_path_wires\[16\]\[7\] VGND VGND VPWR VPWR _02003_
+ sky130_fd_sc_hd__clkbuf_4
Xhold434 top_inst.axis_in_inst.inbuf_bus\[5\] VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1098 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold445 top_inst.deskew_buff_inst.col_input\[109\] VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21181_ _02914_ _02915_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__or2b_1
XFILLER_0_106_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold456 _00964_ VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold467 _00060_ VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap175 net176 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_229_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20132_ _01942_ _01943_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__or2_1
Xhold478 _01165_ VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold489 _00062_ VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_217_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20063_ _01870_ _01877_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_176_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23822_ clknet_leaf_93_clk _00355_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20965_ _02716_ _02732_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__nand2_1
X_23753_ clknet_leaf_122_clk net322 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22704_ _04365_ _04367_ _04376_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_166_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20896_ _02473_ _02646_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__nand2_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23684_ clknet_leaf_117_clk net436 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22635_ _04309_ _04310_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__and2_2
XFILLER_0_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22566_ _04240_ _04244_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__xor2_2
XFILLER_0_10_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24305_ clknet_leaf_2_clk _00838_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[80\]
+ sky130_fd_sc_hd__dfxtp_1
X_21517_ _03244_ _03248_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22497_ _04177_ _04178_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12250_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[15\] _05156_
+ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__or2_1
X_21448_ _03180_ _03182_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__xnor2_2
X_24236_ clknet_leaf_113_clk _00769_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_224_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24167_ clknet_leaf_8_clk _00700_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12181_ top_inst.axis_out_inst.out_buff_data\[18\] _05115_ VGND VGND VPWR VPWR _05118_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_181_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21379_ _03109_ _03111_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23118_ net988 _04656_ _04660_ _04643_ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__o211a_1
X_24098_ clknet_leaf_97_clk _00631_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23049_ net995 _04616_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__or2_1
XTAP_5210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15940_ _08512_ _08513_ _08550_ VGND VGND VPWR VPWR _08551_ sky130_fd_sc_hd__o21a_1
XTAP_5221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15871_ _08444_ _08482_ VGND VGND VPWR VPWR _08483_ sky130_fd_sc_hd__nor2_2
XTAP_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ _10121_ _10122_ VGND VGND VPWR VPWR _10123_ sky130_fd_sc_hd__nor2_1
XFILLER_0_235_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14822_ _07492_ _07507_ VGND VGND VPWR VPWR _07508_ sky130_fd_sc_hd__xnor2_1
XTAP_5298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ _11044_ _11048_ VGND VGND VPWR VPWR _11050_ sky130_fd_sc_hd__or2_1
XTAP_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _10059_ sky130_fd_sc_hd__clkbuf_4
X_14753_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[11\] _07048_ _07438_
+ _07440_ _06180_ VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__o221a_1
XTAP_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ _04994_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13704_ _06417_ _06422_ _06448_ VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__o21a_1
X_17472_ _09998_ _10007_ VGND VGND VPWR VPWR _10008_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_1412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14684_ _07332_ _07340_ VGND VGND VPWR VPWR _07373_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11896_ net670 _04951_ _04954_ _04955_ VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19211_ _11387_ _11590_ _11626_ VGND VGND VPWR VPWR _11627_ sky130_fd_sc_hd__o21a_1
XFILLER_0_157_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16423_ _08984_ _08985_ VGND VGND VPWR VPWR _09002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13635_ _06296_ _06332_ _06381_ VGND VGND VPWR VPWR _06382_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_184_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19142_ _11351_ top_inst.grid_inst.data_path_wires\[13\]\[6\] _11558_ VGND VGND VPWR
+ VPWR _11560_ sky130_fd_sc_hd__o21ai_1
X_16354_ _08882_ VGND VGND VPWR VPWR _08935_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13566_ _06290_ _06291_ _06314_ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_15_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1042 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15305_ _07930_ _07932_ VGND VGND VPWR VPWR _07950_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12517_ _05284_ _05272_ _05332_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__and3_1
X_19073_ _11435_ _11451_ _11450_ VGND VGND VPWR VPWR _11493_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_152_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16285_ _08866_ _08867_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[7\]
+ _07816_ VGND VGND VPWR VPWR _08868_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_70_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13497_ _06245_ _06246_ _06230_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18024_ _10413_ _10524_ VGND VGND VPWR VPWR _10526_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15236_ _07876_ _07882_ VGND VGND VPWR VPWR _07883_ sky130_fd_sc_hd__xor2_1
XFILLER_0_164_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12448_ _05274_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15167_ _05326_ VGND VGND VPWR VPWR _07816_ sky130_fd_sc_hd__buf_6
XFILLER_0_140_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12379_ net418 _05222_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__or2_1
XFILLER_0_205_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14118_ _06823_ _06832_ VGND VGND VPWR VPWR _06833_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_201_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19975_ _01759_ _01758_ _01774_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__a21boi_1
X_15098_ top_inst.grid_inst.data_path_wires\[6\]\[2\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[6\]\[3\]
+ VGND VGND VPWR VPWR _07748_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_240_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14049_ _06762_ _06763_ _06764_ VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__o21a_1
X_18926_ _11161_ _11138_ VGND VGND VPWR VPWR _11349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18857_ _11270_ _11281_ VGND VGND VPWR VPWR _11282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17808_ _10231_ _10261_ _10315_ VGND VGND VPWR VPWR _10316_ sky130_fd_sc_hd__a21oi_1
X_18788_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[3\] _11195_ _11196_
+ VGND VGND VPWR VPWR _11215_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_59_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17739_ _10246_ _10059_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[6\]
+ top_inst.grid_inst.data_path_wires\[11\]\[2\] VGND VGND VPWR VPWR _10248_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_1211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20750_ _02517_ _02519_ _02526_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__a21o_1
XFILLER_0_203_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19409_ _01236_ _01237_ _01244_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20681_ _02365_ _02440_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22420_ _03695_ _03709_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__nand2_2
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22351_ _04034_ _04036_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21302_ _03038_ _03039_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22282_ _03933_ _03934_ _03968_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__and3_1
XFILLER_0_198_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24021_ clknet_leaf_55_clk _00554_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold220 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[6\] VGND
+ VGND VPWR VPWR net402 sky130_fd_sc_hd__dlygate4sd3_1
X_21233_ _02866_ _02887_ _02952_ _02925_ _02891_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__a32o_1
Xhold231 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[3\] VGND VGND
+ VPWR VPWR net413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold242 top_inst.deskew_buff_inst.col_input\[101\] VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold253 top_inst.deskew_buff_inst.col_input\[18\] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _00143_ VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__dlygate4sd3_1
X_21164_ _02906_ _02907_ _05732_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold275 _00266_ VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold286 top_inst.axis_out_inst.out_buff_data\[77\] VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 _00074_ VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_244_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20115_ _01903_ _01926_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21095_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[31\] _02856_ VGND
+ VGND VPWR VPWR _02857_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_244_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20046_ _01841_ _01842_ _01860_ _10957_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__a31o_1
XFILLER_0_217_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23805_ clknet_leaf_69_clk _00338_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 _05275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_217_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_1418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_115 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ _03700_ _05275_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__or2_1
XFILLER_0_233_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ net451 _04865_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__or2_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23736_ clknet_leaf_125_clk _00269_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ _02643_ _02693_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23667_ clknet_leaf_124_clk _00200_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20879_ _02528_ _02644_ _02650_ VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__a21o_1
XFILLER_0_193_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13420_ top_inst.grid_inst.data_path_wires\[2\]\[3\] VGND VGND VPWR VPWR _06188_
+ sky130_fd_sc_hd__buf_4
XFILLER_0_14_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22618_ _04287_ _04294_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23598_ clknet_leaf_101_clk _00131_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13351_ _06123_ _06124_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22549_ _04203_ _04191_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12302_ net874 _05178_ _05187_ _05182_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__o211a_1
XFILLER_0_228_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16070_ _08671_ _08140_ VGND VGND VPWR VPWR _08672_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13282_ _06013_ _06014_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__or2b_1
XFILLER_0_133_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15021_ _07613_ _07610_ _07629_ _07627_ VGND VGND VPWR VPWR _07674_ sky130_fd_sc_hd__nand4_1
X_24219_ clknet_leaf_19_clk _00752_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12233_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[8\] _05143_
+ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12164_ top_inst.axis_out_inst.out_buff_data\[11\] _05102_ VGND VGND VPWR VPWR _05108_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_31_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16972_ _09499_ _09525_ _09526_ VGND VGND VPWR VPWR _09527_ sky130_fd_sc_hd__and3_1
X_19760_ _01565_ _01587_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__xnor2_2
X_12095_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[13\] _05063_
+ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__or2_1
XFILLER_0_235_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18711_ _05772_ VGND VGND VPWR VPWR _11150_ sky130_fd_sc_hd__clkbuf_4
X_15923_ _08532_ _08533_ VGND VGND VPWR VPWR _08534_ sky130_fd_sc_hd__nor2_1
XTAP_5040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19691_ _01476_ _01505_ _01504_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_127_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18642_ _11098_ _11052_ VGND VGND VPWR VPWR _11100_ sky130_fd_sc_hd__nand2_1
XTAP_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _08429_ _08466_ VGND VGND VPWR VPWR _08467_ sky130_fd_sc_hd__and2_1
XTAP_5095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_203_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14805_ _07489_ _07490_ VGND VGND VPWR VPWR _07491_ sky130_fd_sc_hd__nor2_1
XTAP_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ _11031_ _11032_ VGND VGND VPWR VPWR _11034_ sky130_fd_sc_hd__nand2_1
XTAP_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15785_ top_inst.grid_inst.data_path_wires\[7\]\[3\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[6\]
+ _08353_ top_inst.grid_inst.data_path_wires\[7\]\[2\] VGND VGND VPWR VPWR _08399_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_207_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12997_ _05738_ _05759_ _05775_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__and3_1
XFILLER_0_231_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17524_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _10047_ sky130_fd_sc_hd__clkbuf_4
XTAP_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_231_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14736_ _07415_ _07423_ VGND VGND VPWR VPWR _07424_ sky130_fd_sc_hd__xnor2_1
XTAP_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11948_ net731 _04982_ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17455_ net1030 _08183_ _09991_ _09231_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__o211a_1
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ _07314_ _07355_ _07057_ VGND VGND VPWR VPWR _07357_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11879_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[16\] _04943_
+ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__or2_1
X_16406_ _08984_ _08985_ VGND VGND VPWR VPWR _08986_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_223_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13618_ _06357_ _06355_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__or2b_1
X_17386_ _09910_ _09925_ VGND VGND VPWR VPWR _09926_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_172_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14598_ _07285_ _07288_ VGND VGND VPWR VPWR _07289_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_82_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19125_ _11505_ _11543_ VGND VGND VPWR VPWR _11544_ sky130_fd_sc_hd__nand2_1
X_16337_ _08870_ _08917_ _08918_ _08692_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13549_ top_inst.grid_inst.data_path_wires\[2\]\[2\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[2\]\[3\]
+ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19056_ _11470_ _11475_ VGND VGND VPWR VPWR _11476_ sky130_fd_sc_hd__xnor2_1
X_16268_ _08801_ _08803_ _08849_ _08850_ VGND VGND VPWR VPWR _08851_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_70_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18007_ _10508_ _10509_ VGND VGND VPWR VPWR _10510_ sky130_fd_sc_hd__nand2_1
XFILLER_0_207_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15219_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[8\] _07866_ VGND
+ VGND VPWR VPWR _07867_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16199_ _08755_ _08757_ VGND VGND VPWR VPWR _08784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_239_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19958_ net1095 _01202_ _01776_ _01777_ _11228_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__o221a_1
X_18909_ _10641_ _11332_ VGND VGND VPWR VPWR _11333_ sky130_fd_sc_hd__and2_1
XFILLER_0_208_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19889_ _01709_ _01711_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_241_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21920_ _03635_ _03636_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21851_ _03549_ _03568_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20802_ _02574_ _02575_ _02465_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24570_ clknet_leaf_134_clk _01103_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dfxtp_2
X_21782_ _03481_ _03505_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23521_ clknet_leaf_139_clk net545 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20733_ _02494_ _02510_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_148_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23452_ net923 _04840_ _04848_ _04844_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20664_ _02426_ _02427_ _02443_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_1337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22403_ net659 _09804_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23383_ net725 _04804_ _04811_ _04808_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__o211a_1
X_20595_ _02374_ _02376_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22334_ _04016_ _04019_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22265_ top_inst.grid_inst.data_path_wires\[18\]\[2\] _03713_ VGND VGND VPWR VPWR
+ _03953_ sky130_fd_sc_hd__and2b_1
XFILLER_0_60_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24004_ clknet_leaf_82_clk _00537_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_131_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21216_ _02932_ _02933_ _02956_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_108_1277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22196_ _03885_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_1422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21147_ _02873_ _02881_ _02894_ _02880_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__o211a_1
XFILLER_0_217_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21078_ _02674_ _02789_ _02786_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_233_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12920_ _05722_ _05723_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__xnor2_1
X_20029_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[24\] _01761_ _01762_
+ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12851_ _05657_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_198_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11802_ _04874_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__clkbuf_4
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _08189_ _08190_ VGND VGND VPWR VPWR _08191_ sky130_fd_sc_hd__or2_1
X_12782_ _05562_ _05554_ _05590_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__a21oi_2
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _07211_ _07212_ _07178_ VGND VGND VPWR VPWR _07214_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_185_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11733_ net35 net166 VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__nor2b_4
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23719_ clknet_leaf_120_clk _00252_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17240_ _09786_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[4\] _07060_ _07064_
+ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _07147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13403_ _06173_ _06174_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17171_ _09698_ _09696_ _09714_ VGND VGND VPWR VPWR _09720_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14383_ _05290_ _07082_ _07084_ _06684_ VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16122_ _08688_ _08661_ VGND VGND VPWR VPWR _08710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13334_ _06080_ _06077_ _06108_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16053_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[16\] _07866_ VGND
+ VGND VPWR VPWR _08660_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13265_ _06041_ VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15004_ _07656_ _07657_ VGND VGND VPWR VPWR _07658_ sky130_fd_sc_hd__nand2_1
X_12216_ net642 _05129_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13196_ _05972_ _05973_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19812_ _01606_ _01609_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12147_ net750 _05097_ _05098_ _05088_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19743_ _01298_ _01314_ _11704_ _11708_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__or4b_1
X_16955_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[5\] _09209_ VGND
+ VGND VPWR VPWR _09510_ sky130_fd_sc_hd__and2_1
X_12078_ net797 _05058_ _05059_ _05049_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15906_ _08152_ _08167_ VGND VGND VPWR VPWR _08517_ sky130_fd_sc_hd__nand2_2
X_16886_ _09386_ _09388_ _09441_ _09442_ VGND VGND VPWR VPWR _09443_ sky130_fd_sc_hd__a211oi_2
X_19674_ _01456_ _01477_ _01502_ _01503_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15837_ _08448_ _08436_ VGND VGND VPWR VPWR _08450_ sky130_fd_sc_hd__and2b_1
X_18625_ _11082_ _11083_ VGND VGND VPWR VPWR _11084_ sky130_fd_sc_hd__or2_1
XTAP_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15768_ _08310_ _08322_ VGND VGND VPWR VPWR _08383_ sky130_fd_sc_hd__nand2_1
X_18556_ _10975_ _11016_ VGND VGND VPWR VPWR _11017_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_172_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14719_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[11\] _07281_ VGND
+ VGND VPWR VPWR _07407_ sky130_fd_sc_hd__xnor2_1
X_17507_ top_inst.grid_inst.data_path_wires\[11\]\[5\] VGND VGND VPWR VPWR _10035_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18487_ _10909_ _10884_ VGND VGND VPWR VPWR _10950_ sky130_fd_sc_hd__or2b_1
XFILLER_0_185_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15699_ _08313_ _08314_ VGND VGND VPWR VPWR _08315_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17438_ _09915_ _09973_ VGND VGND VPWR VPWR _09975_ sky130_fd_sc_hd__nand2_1
XANTENNA_15 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_26 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_37 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_48 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17369_ _09892_ _09905_ VGND VGND VPWR VPWR _09909_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_59 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19108_ _11480_ _11482_ VGND VGND VPWR VPWR _11527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20380_ _02164_ _02165_ _02104_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_207_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19039_ _11420_ _11459_ VGND VGND VPWR VPWR _11460_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput100 net100 VGND VGND VPWR VPWR output_tdata[40] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput111 net111 VGND VGND VPWR VPWR output_tdata[50] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput122 net122 VGND VGND VPWR VPWR output_tdata[60] sky130_fd_sc_hd__buf_2
Xoutput133 net133 VGND VGND VPWR VPWR output_tdata[70] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22050_ _03686_ _03684_ _03700_ _03698_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__nand4_1
XFILLER_0_140_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput144 net144 VGND VGND VPWR VPWR output_tdata[80] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput155 net155 VGND VGND VPWR VPWR output_tdata[90] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput166 net166 VGND VGND VPWR VPWR output_tvalid sky130_fd_sc_hd__clkbuf_4
X_21001_ _02463_ _02747_ _02503_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22952_ net416 _04557_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21903_ _03453_ _03581_ _03598_ _03601_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__o31a_1
XFILLER_0_218_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22883_ net294 _04522_ _04525_ _04524_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24622_ clknet_leaf_22_clk net532 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[98\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21834_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[23\] _03421_ _03422_
+ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_210_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24553_ clknet_leaf_103_clk _01086_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_78_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21765_ net886 _06169_ _03489_ _02909_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23504_ clknet_leaf_139_clk _00037_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[94\]
+ sky130_fd_sc_hd__dfxtp_2
X_20716_ _02484_ _02483_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__or2b_1
XFILLER_0_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24484_ clknet_leaf_115_clk _01017_ VGND VGND VPWR VPWR top_inst.valid_pipe\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21696_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[17\] _03421_ _03422_
+ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_108_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23435_ net443 _04835_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20647_ _02403_ _02410_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_983 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23366_ net444 _04791_ _04801_ _04795_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__o211a_1
X_20578_ _01997_ _02229_ _02357_ _02358_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__nor4_1
XFILLER_0_190_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22317_ _03976_ _04003_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__xnor2_2
X_23297_ net468 _04752_ _04762_ _04756_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__o211a_1
XFILLER_0_225_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13050_ top_inst.grid_inst.data_path_wires\[1\]\[5\] top_inst.grid_inst.data_path_wires\[1\]\[4\]
+ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__and4_1
XFILLER_0_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22248_ _03890_ _03895_ _03935_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12001_ net497 _05004_ _05015_ _05008_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__o211a_1
X_22179_ _03867_ _03868_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16740_ _09268_ _09270_ _09298_ _09299_ VGND VGND VPWR VPWR _09300_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13952_ top_inst.grid_inst.data_path_wires\[3\]\[3\] top_inst.grid_inst.data_path_wires\[3\]\[2\]
+ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _06672_ sky130_fd_sc_hd__and4_1
XFILLER_0_57_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12903_ _05706_ _05707_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__and2_1
XFILLER_0_199_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_214_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16671_ _09194_ _09189_ _09192_ _09197_ VGND VGND VPWR VPWR _09234_ sky130_fd_sc_hd__nand4_2
XFILLER_0_220_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13883_ _06181_ _06192_ _06621_ _06446_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__o211a_1
XFILLER_0_232_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18410_ _10871_ _10873_ VGND VGND VPWR VPWR _10875_ sky130_fd_sc_hd__and2_1
X_15622_ top_inst.grid_inst.data_path_wires\[7\]\[1\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[7\]\[2\]
+ VGND VGND VPWR VPWR _08240_ sky130_fd_sc_hd__a22o_1
X_12834_ top_inst.axis_in_inst.inbuf_bus\[6\] _05267_ _05640_ VGND VGND VPWR VPWR
+ _05641_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19390_ net355 _01202_ _01225_ _01226_ _11228_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__o221a_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _10599_ _10612_ _10769_ VGND VGND VPWR VPWR _10807_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15553_ _08135_ _08157_ _08155_ _08137_ VGND VGND VPWR VPWR _08175_ sky130_fd_sc_hd__a22o_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _05293_ _05301_ _05306_ _05288_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_201_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14504_ _07194_ _07195_ _07172_ _07173_ VGND VGND VPWR VPWR _07197_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_167_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18272_ _10737_ _10738_ _10713_ _10714_ VGND VGND VPWR VPWR _10740_ sky130_fd_sc_hd__o211a_1
X_15484_ _08110_ _08111_ _08123_ VGND VGND VPWR VPWR _08124_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12696_ _05280_ _05273_ _05305_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17223_ _09752_ _09757_ _09755_ VGND VGND VPWR VPWR _09770_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_182_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14435_ _07118_ _07111_ _07129_ VGND VGND VPWR VPWR _07131_ sky130_fd_sc_hd__or3_1
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput13 input_tdata[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17154_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[15\] _09631_ VGND
+ VGND VPWR VPWR _09704_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput24 input_tdata[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14366_ _07070_ _06641_ VGND VGND VPWR VPWR _07071_ sky130_fd_sc_hd__or2_1
Xinput35 output_tready VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_4
XFILLER_0_107_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_208_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16105_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _08697_ sky130_fd_sc_hd__buf_2
X_13317_ _06054_ _06091_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__xnor2_1
Xhold808 top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[0\] VGND VGND
+ VPWR VPWR net990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17085_ _09361_ _09215_ _09219_ _09213_ VGND VGND VPWR VPWR _09637_ sky130_fd_sc_hd__a2bb2o_1
Xhold819 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[1\] VGND
+ VGND VPWR VPWR net1001 sky130_fd_sc_hd__dlygate4sd3_1
X_14297_ _07005_ _07006_ VGND VGND VPWR VPWR _07007_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16036_ _08614_ _08616_ _08643_ VGND VGND VPWR VPWR _08644_ sky130_fd_sc_hd__o21ba_1
X_13248_ _05945_ _06024_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__nor2_1
XFILLER_0_228_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13179_ _05865_ _05909_ _05957_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_237_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17987_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[13\] _10367_ _10283_
+ VGND VGND VPWR VPWR _10490_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19726_ _01519_ _01553_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16938_ _05312_ VGND VGND VPWR VPWR _09494_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_237_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19657_ _01484_ _01485_ _01402_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__o21ai_4
X_16869_ _09424_ _09425_ VGND VGND VPWR VPWR _09426_ sky130_fd_sc_hd__nor2_1
XFILLER_0_232_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18608_ _11027_ _11066_ _11067_ VGND VGND VPWR VPWR _11068_ sky130_fd_sc_hd__a21oi_2
X_19588_ net249 _01418_ _01419_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__and3_1
XFILLER_0_181_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18539_ _10999_ _11000_ VGND VGND VPWR VPWR _11001_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21550_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[13\] _03080_ VGND
+ VGND VPWR VPWR _03282_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_691 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20501_ _01997_ _02018_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21481_ _03211_ _03214_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23220_ net610 _04713_ _04719_ _04717_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__o211a_1
X_20432_ _02176_ _02217_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_244_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23151_ net72 _04672_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__or2_1
X_20363_ top_inst.grid_inst.data_path_wires\[16\]\[3\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[3\]
+ _02051_ top_inst.grid_inst.data_path_wires\[16\]\[4\] VGND VGND VPWR VPWR _02150_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22102_ _03785_ _03793_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__xor2_2
X_23082_ top_inst.axis_in_inst.inbuf_bus\[28\] _04629_ VGND VGND VPWR VPWR _04639_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_113_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20294_ _02077_ _02054_ _02081_ _02082_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22033_ _03726_ _03727_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__nand2_1
XTAP_6329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23984_ clknet_leaf_80_clk _00517_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_242_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1056 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22935_ net612 _04543_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__or2_1
XFILLER_0_202_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22866_ net1006 _04509_ _04515_ _04511_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24605_ clknet_leaf_21_clk _01138_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_210_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21817_ _03537_ _03538_ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_1380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22797_ net564 _06169_ _04465_ _03929_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12550_ _05363_ _05284_ _05283_ _05364_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__and4b_1
X_24536_ clknet_leaf_102_clk _01069_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dfxtp_2
XPHY_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21748_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[19\] _03421_ _03422_
+ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__a21oi_2
XPHY_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24467_ clknet_leaf_55_clk _01000_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_12481_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _05302_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21679_ _03246_ _03406_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14220_ _06930_ _06931_ VGND VGND VPWR VPWR _06932_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23418_ net531 _04827_ _04829_ _04819_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24398_ clknet_leaf_38_clk _00931_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_1113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14151_ _06811_ _06863_ _06864_ VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_34_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23349_ _04686_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__buf_2
XFILLER_0_22_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13102_ _05325_ _05882_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14082_ _06795_ _06797_ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_162_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_219_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13033_ _05802_ _05815_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__xnor2_1
X_17910_ _10413_ _10414_ VGND VGND VPWR VPWR _10415_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18890_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[5\] _11135_ VGND
+ VGND VPWR VPWR _11314_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17841_ _10333_ _10334_ _10346_ VGND VGND VPWR VPWR _10348_ sky130_fd_sc_hd__and3_1
XFILLER_0_234_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17772_ _10237_ _10233_ VGND VGND VPWR VPWR _10280_ sky130_fd_sc_hd__or2b_1
X_14984_ _07640_ _07641_ VGND VGND VPWR VPWR _07642_ sky130_fd_sc_hd__or2_1
XFILLER_0_234_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19511_ _01344_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__clkbuf_1
X_16723_ _09256_ VGND VGND VPWR VPWR _09284_ sky130_fd_sc_hd__inv_2
X_13935_ _06622_ _06637_ _06618_ _06640_ VGND VGND VPWR VPWR _06657_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16654_ _05269_ _09219_ VGND VGND VPWR VPWR _09220_ sky130_fd_sc_hd__or2_1
XFILLER_0_159_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19442_ _01272_ _01273_ _01276_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__nand3_1
X_13866_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[14\] _06242_ _06605_
+ _06606_ VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15605_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[3\] _08203_ _08204_
+ VGND VGND VPWR VPWR _08224_ sky130_fd_sc_hd__a21bo_1
X_12817_ _05582_ _05623_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16585_ _09126_ _09129_ _09128_ VGND VGND VPWR VPWR _09160_ sky130_fd_sc_hd__o21ba_1
X_19373_ _01207_ _01208_ _01209_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__nand3_1
XFILLER_0_9_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13797_ _06538_ _06458_ net181 VGND VGND VPWR VPWR _06540_ sky130_fd_sc_hd__or3_2
XFILLER_0_158_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18324_ _10763_ _10765_ VGND VGND VPWR VPWR _10790_ sky130_fd_sc_hd__nand2_1
X_15536_ top_inst.grid_inst.data_path_wires\[7\]\[4\] VGND VGND VPWR VPWR _08163_
+ sky130_fd_sc_hd__buf_4
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12748_ _05520_ _05522_ _05556_ _05557_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_31_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18255_ _10716_ _10722_ VGND VGND VPWR VPWR _10723_ sky130_fd_sc_hd__xnor2_1
X_15467_ _08102_ _08106_ VGND VGND VPWR VPWR _08108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_210_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12679_ _05282_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17206_ _09588_ _09459_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[17\]
+ VGND VGND VPWR VPWR _09754_ sky130_fd_sc_hd__a21o_1
XFILLER_0_170_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14418_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[2\] _06242_ _07113_
+ _07114_ VGND VGND VPWR VPWR _07115_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18186_ _10656_ VGND VGND VPWR VPWR _10657_ sky130_fd_sc_hd__inv_2
X_15398_ _08030_ _07998_ _08040_ VGND VGND VPWR VPWR _08041_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17137_ _09686_ _09687_ VGND VGND VPWR VPWR _09688_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14349_ _05731_ VGND VGND VPWR VPWR _07057_ sky130_fd_sc_hd__buf_8
XFILLER_0_25_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold605 top_inst.axis_out_inst.out_buff_data\[1\] VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 _00140_ VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold627 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[4\] VGND VGND
+ VPWR VPWR net809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold638 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[30\] VGND
+ VGND VPWR VPWR net820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17068_ _08870_ _09619_ _09620_ _09231_ VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__o211a_1
Xhold649 top_inst.axis_out_inst.out_buff_data\[93\] VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16019_ _08601_ _08608_ _08600_ VGND VGND VPWR VPWR _08627_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19709_ _01535_ _01536_ _01534_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_1365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20981_ _02528_ _02741_ _02748_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_240_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22720_ _04390_ _04391_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22651_ _04284_ _04301_ _04322_ _04325_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_149_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21602_ _03284_ _03285_ _03298_ _03297_ _03295_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__o32a_1
X_22582_ _04256_ _04253_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__or2b_1
XFILLER_0_76_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24321_ clknet_leaf_9_clk _00854_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[18\]\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_21533_ _03205_ _03206_ _03222_ _03221_ _03219_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__o32a_1
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24252_ clknet_leaf_107_clk _00785_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21464_ _03188_ _03161_ VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__or2b_1
XFILLER_0_181_1216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23203_ net378 _04700_ _04709_ _04704_ VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20415_ _02148_ _02156_ _02155_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_209_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24183_ clknet_leaf_29_clk _00716_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21395_ top_inst.grid_inst.data_path_wires\[17\]\[5\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[17\]\[6\]
+ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_226_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23134_ net154 _04659_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20346_ top_inst.deskew_buff_inst.col_input\[37\] _05634_ _02132_ _02133_ VGND VGND
+ VPWR VPWR _02134_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_102_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23065_ net590 _04629_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__or2_1
X_20277_ _02063_ _02064_ _02065_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__a21oi_1
XTAP_6126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22016_ _03713_ _05275_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__or2_1
XFILLER_0_234_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_236_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23967_ clknet_leaf_90_clk _00500_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_11981_ net551 _04990_ _05003_ _04995_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_242_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13720_ _06463_ _06464_ VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__nor2_1
X_22918_ top_inst.skew_buff_inst.row\[2\].output_reg\[6\] _04543_ VGND VGND VPWR VPWR
+ _04545_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23898_ clknet_leaf_52_clk _00431_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13651_ _06306_ _06348_ _06397_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__a21boi_1
X_22849_ net715 _04504_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__or2_1
XFILLER_0_211_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12602_ _05413_ _05414_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16370_ _08908_ _08909_ _08950_ VGND VGND VPWR VPWR _08951_ sky130_fd_sc_hd__o21a_1
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_1097 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13582_ _06328_ _06329_ VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15321_ _07956_ _07964_ VGND VGND VPWR VPWR _07966_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12533_ _05347_ _05348_ VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__nor2_1
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24519_ clknet_leaf_132_clk _01052_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_152_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18040_ _10520_ _10539_ _10540_ _10541_ _04861_ VGND VGND VPWR VPWR _10542_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_227_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15252_ _07853_ _07855_ VGND VGND VPWR VPWR _07899_ sky130_fd_sc_hd__or2_1
X_12464_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _05288_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_163_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14203_ _06875_ _06877_ _06915_ VGND VGND VPWR VPWR _06916_ sky130_fd_sc_hd__o21a_1
XFILLER_0_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15183_ _07828_ _07830_ VGND VGND VPWR VPWR _07831_ sky130_fd_sc_hd__xnor2_2
X_12395_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[14\] _05235_
+ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14134_ _05732_ VGND VGND VPWR VPWR _06848_ sky130_fd_sc_hd__buf_4
X_19991_ _01800_ _01808_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14065_ _06775_ _06780_ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__xnor2_2
X_18942_ _11362_ _11364_ VGND VGND VPWR VPWR _11365_ sky130_fd_sc_hd__xor2_1
XFILLER_0_123_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13016_ _05785_ _05798_ _05797_ VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__o21a_1
XFILLER_0_197_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18873_ _11263_ _11269_ VGND VGND VPWR VPWR _11297_ sky130_fd_sc_hd__or2b_1
XFILLER_0_123_1199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17824_ _10329_ _10330_ VGND VGND VPWR VPWR _10331_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14967_ _07629_ _07075_ VGND VGND VPWR VPWR _07630_ sky130_fd_sc_hd__or2_1
X_17755_ _10219_ _10194_ VGND VGND VPWR VPWR _10264_ sky130_fd_sc_hd__or2b_1
XFILLER_0_206_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16706_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[2\] _09197_ VGND
+ VGND VPWR VPWR _09267_ sky130_fd_sc_hd__nand2_1
X_13918_ _06645_ _06641_ VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__or2_1
X_14898_ _07450_ _07562_ _07580_ VGND VGND VPWR VPWR _07581_ sky130_fd_sc_hd__o21ai_1
X_17686_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[6\] _10161_ _10162_
+ VGND VGND VPWR VPWR _10196_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19425_ _01247_ _01248_ _01249_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__nor3b_1
X_16637_ net216 VGND VGND VPWR VPWR _09206_ sky130_fd_sc_hd__buf_4
X_13849_ _06198_ _06524_ _06527_ _06557_ VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_230_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_943 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19356_ _01186_ _01193_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16568_ _09066_ _09068_ _09110_ _09111_ _09113_ VGND VGND VPWR VPWR _09144_ sky130_fd_sc_hd__a32o_1
XFILLER_0_146_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18307_ _10761_ _10773_ VGND VGND VPWR VPWR _10774_ sky130_fd_sc_hd__xnor2_1
X_15519_ _07622_ _06634_ _08151_ _08142_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16499_ _09075_ _09076_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[12\]
+ _07816_ VGND VGND VPWR VPWR _09077_ sky130_fd_sc_hd__a2bb2o_1
X_19287_ _05772_ VGND VGND VPWR VPWR _11689_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_161_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18238_ _10682_ _10706_ VGND VGND VPWR VPWR _10707_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18169_ _10071_ _10638_ _10640_ _10620_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__o211a_1
Xhold402 _00972_ VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold413 top_inst.axis_out_inst.out_buff_data\[40\] VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__dlygate4sd3_1
X_20200_ _02001_ _05739_ _02002_ _01840_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__o211a_1
Xhold424 top_inst.axis_in_inst.inbuf_bus\[8\] VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__dlygate4sd3_1
X_21180_ _02907_ _02919_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__or2b_1
Xhold435 _00979_ VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold446 _01166_ VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold457 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[24\] VGND VGND
+ VPWR VPWR net639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20131_ _01918_ _01933_ _01941_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__and3_1
Xhold468 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[22\] VGND
+ VGND VPWR VPWR net650 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap176 _02320_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold479 top_inst.axis_out_inst.out_buff_data\[9\] VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20062_ _01876_ _01868_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__xor2_2
XFILLER_0_96_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_225_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23821_ clknet_leaf_93_clk _00354_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23752_ clknet_leaf_122_clk net334 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20964_ _02716_ _02732_ VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__or2_2
XFILLER_0_67_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22703_ _04368_ _04375_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__xnor2_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23683_ clknet_leaf_119_clk _00216_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20895_ _02466_ _02468_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22634_ _04218_ _04308_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22565_ _04242_ _04243_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24304_ clknet_leaf_2_clk _00837_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[79\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_1081 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21516_ _03244_ _03248_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__and2_1
XFILLER_0_161_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22496_ _04174_ _04176_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__and2_1
XFILLER_0_161_642 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24235_ clknet_leaf_113_clk _00768_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_21447_ _03136_ _03144_ _03181_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_181_1035 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24166_ clknet_leaf_9_clk _00699_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[8\]
+ sky130_fd_sc_hd__dfxtp_2
X_12180_ net885 _05110_ _05117_ _05114_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__o211a_1
X_21378_ _03070_ _03113_ _03114_ _02909_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23117_ net38 _04659_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__or2_1
X_20329_ _02108_ _02115_ _02116_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__nand3_1
X_24097_ clknet_leaf_99_clk _00630_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23048_ net4 _04615_ _04620_ _04619_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__o211a_1
XTAP_5200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15870_ _08164_ _08161_ top_inst.grid_inst.data_path_wires\[7\]\[7\] VGND VGND VPWR
+ VPWR _08482_ sky130_fd_sc_hd__o21ai_1
XTAP_5255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14821_ _07505_ _07506_ VGND VGND VPWR VPWR _07507_ sky130_fd_sc_hd__nand2_1
XFILLER_0_216_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_243_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14752_ _07398_ _07403_ net1124 _07439_ VGND VGND VPWR VPWR _07440_ sky130_fd_sc_hd__a31o_1
XTAP_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17540_ _10038_ _10046_ _10058_ _10049_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__o211a_1
XTAP_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _04873_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _06416_ _06415_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__or2b_1
XFILLER_0_86_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17471_ _10005_ _10006_ VGND VGND VPWR VPWR _10007_ sky130_fd_sc_hd__and2_1
XTAP_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14683_ _07338_ _07339_ VGND VGND VPWR VPWR _07372_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_230_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11895_ _04874_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_1424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19210_ _11624_ _11625_ VGND VGND VPWR VPWR _11626_ sky130_fd_sc_hd__nor2_1
X_16422_ _08981_ _08983_ VGND VGND VPWR VPWR _09001_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13634_ _06333_ _06336_ _06337_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16353_ _08927_ _08933_ VGND VGND VPWR VPWR _08934_ sky130_fd_sc_hd__xor2_1
X_19141_ _11351_ top_inst.grid_inst.data_path_wires\[13\]\[6\] _11558_ VGND VGND VPWR
+ VPWR _11559_ sky130_fd_sc_hd__or3_1
XFILLER_0_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13565_ _06293_ _06313_ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__xor2_1
XFILLER_0_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15304_ _07935_ _07937_ VGND VGND VPWR VPWR _07949_ sky130_fd_sc_hd__nor2_1
X_12516_ _05284_ _05272_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__a21oi_1
X_19072_ _11476_ _11491_ VGND VGND VPWR VPWR _11492_ sky130_fd_sc_hd__xor2_1
X_16284_ _08864_ _08865_ _05353_ VGND VGND VPWR VPWR _08867_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13496_ _06230_ _06245_ _06246_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15235_ _07880_ _07881_ VGND VGND VPWR VPWR _07882_ sky130_fd_sc_hd__xor2_1
X_18023_ _10413_ _10524_ VGND VGND VPWR VPWR _10525_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12447_ top_inst.axis_in_inst.inbuf_valid _05267_ _04857_ VGND VGND VPWR VPWR _05274_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_129_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15166_ _07812_ _07813_ _06404_ VGND VGND VPWR VPWR _07815_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12378_ _05177_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__buf_2
XFILLER_0_205_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14117_ _06829_ _06831_ VGND VGND VPWR VPWR _06832_ sky130_fd_sc_hd__nor2_1
X_19974_ _01749_ _01775_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__and2_1
X_15097_ _07745_ _07746_ VGND VGND VPWR VPWR _07747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14048_ _06762_ _06763_ _06764_ VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__nor3_1
X_18925_ _11346_ _11347_ VGND VGND VPWR VPWR _11348_ sky130_fd_sc_hd__nand2_1
XFILLER_0_238_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18856_ _11271_ _11280_ VGND VGND VPWR VPWR _11281_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17807_ _10258_ _10260_ VGND VGND VPWR VPWR _10315_ sky130_fd_sc_hd__nor2_1
XFILLER_0_238_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18787_ _11193_ _11213_ VGND VGND VPWR VPWR _11214_ sky130_fd_sc_hd__xor2_2
XFILLER_0_55_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15999_ _08603_ _08607_ VGND VGND VPWR VPWR _08608_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17738_ top_inst.grid_inst.data_path_wires\[11\]\[2\] _10246_ _10059_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _10247_ sky130_fd_sc_hd__and4_1
XFILLER_0_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17669_ _10158_ _10178_ _10179_ VGND VGND VPWR VPWR _10180_ sky130_fd_sc_hd__and3_1
XFILLER_0_187_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19408_ _01242_ _01243_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20680_ _02428_ _02435_ _02458_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19339_ net172 _11732_ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22350_ _03986_ _03994_ _04035_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_127_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21301_ _02878_ _02875_ _02885_ _02883_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__nand4_1
XFILLER_0_143_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_889 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22281_ _03933_ _03934_ _03968_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24020_ clknet_leaf_54_clk _00553_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_5_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold210 top_inst.axis_out_inst.out_buff_data\[113\] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21232_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[4\] _02944_ _02945_
+ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__a21boi_2
Xhold221 _00173_ VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 _00937_ VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold243 _01158_ VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold254 _00217_ VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[1\] VGND
+ VGND VPWR VPWR net447 sky130_fd_sc_hd__dlygate4sd3_1
X_21163_ _02899_ _02904_ _02905_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__nand3_2
XFILLER_0_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold276 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[6\] VGND
+ VGND VPWR VPWR net458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold287 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[21\] VGND
+ VGND VPWR VPWR net469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20114_ _01903_ _01926_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__nand2_1
Xhold298 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[16\] VGND
+ VGND VPWR VPWR net480 sky130_fd_sc_hd__dlygate4sd3_1
X_21094_ _02854_ _02855_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_244_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_217_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20045_ _01841_ _01842_ _01860_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__a21oi_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23804_ clknet_leaf_77_clk _00337_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 _05275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21996_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _03700_ sky130_fd_sc_hd__clkbuf_4
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23735_ clknet_leaf_126_clk net453 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ _02701_ _02700_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__or2b_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23666_ clknet_leaf_124_clk _00199_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20878_ _02463_ _02649_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22617_ _04293_ _04285_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__xor2_2
XFILLER_0_14_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23597_ clknet_leaf_101_clk _00130_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13350_ _06054_ _06122_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__or2_1
XFILLER_0_181_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22548_ _04202_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12301_ net452 _05183_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13281_ _06055_ _06056_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22479_ _04127_ _04130_ _04129_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15020_ _07610_ _07629_ _07627_ _07613_ VGND VGND VPWR VPWR _07673_ sky130_fd_sc_hd__a22o_1
X_24218_ clknet_leaf_19_clk _00751_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12232_ net585 _05137_ _05147_ _05141_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__o211a_1
XFILLER_0_224_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24149_ clknet_leaf_17_clk _00682_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[13\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12163_ net357 _05097_ _05107_ _05101_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16971_ _09523_ _09524_ _09481_ _09500_ VGND VGND VPWR VPWR _09526_ sky130_fd_sc_hd__o211ai_2
X_12094_ net439 _05058_ _05068_ _05062_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18710_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _11149_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15922_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[12\] _08374_ VGND
+ VGND VPWR VPWR _08533_ sky130_fd_sc_hd__xnor2_1
XTAP_5041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19690_ _01508_ _01509_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__nand2_1
XTAP_5052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18641_ _11098_ _11055_ _11077_ _11084_ VGND VGND VPWR VPWR _11099_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_239_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15853_ _08463_ _08465_ VGND VGND VPWR VPWR _08466_ sky130_fd_sc_hd__xor2_1
XFILLER_0_244_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14804_ _07450_ _07488_ VGND VGND VPWR VPWR _07490_ sky130_fd_sc_hd__and2_1
XTAP_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18572_ _11031_ _11032_ VGND VGND VPWR VPWR _11033_ sky130_fd_sc_hd__or2_1
X_12996_ _05741_ _05757_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__nand2_1
XTAP_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15784_ top_inst.grid_inst.data_path_wires\[7\]\[2\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[7\]
+ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[7\]\[3\]
+ VGND VGND VPWR VPWR _08398_ sky130_fd_sc_hd__and4b_1
XFILLER_0_99_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17523_ _05755_ VGND VGND VPWR VPWR _10046_ sky130_fd_sc_hd__clkbuf_4
XTAP_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14735_ _07421_ _07422_ VGND VGND VPWR VPWR _07423_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11947_ net549 _04977_ _04984_ _04981_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _07314_ _07355_ VGND VGND VPWR VPWR _07356_ sky130_fd_sc_hd__nor2_1
X_17454_ _09984_ _09985_ _09990_ _05732_ VGND VGND VPWR VPWR _09991_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11878_ net544 _04938_ _04945_ _04942_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16405_ _08938_ _08942_ _08940_ VGND VGND VPWR VPWR _08985_ sky130_fd_sc_hd__a21oi_1
X_13617_ _04869_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__buf_4
XFILLER_0_144_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14597_ _07286_ _07287_ VGND VGND VPWR VPWR _07288_ sky130_fd_sc_hd__nor2_1
X_17385_ _09922_ _09924_ VGND VGND VPWR VPWR _09925_ sky130_fd_sc_hd__xor2_1
XFILLER_0_223_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19124_ _11498_ _11542_ VGND VGND VPWR VPWR _11543_ sky130_fd_sc_hd__xnor2_1
X_16336_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[8\] _07866_ VGND
+ VGND VPWR VPWR _08918_ sky130_fd_sc_hd__or2_1
X_13548_ _06295_ _06296_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16267_ _08847_ _08848_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[7\]
+ VGND VGND VPWR VPWR _08850_ sky130_fd_sc_hd__a21oi_1
X_19055_ _11473_ _11474_ VGND VGND VPWR VPWR _11475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_242_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13479_ _06229_ _06230_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__or2_1
XFILLER_0_207_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15218_ _05312_ VGND VGND VPWR VPWR _07866_ sky130_fd_sc_hd__clkbuf_4
X_18006_ _10507_ _10489_ VGND VGND VPWR VPWR _10509_ sky130_fd_sc_hd__or2b_1
X_16198_ _08780_ _08782_ VGND VGND VPWR VPWR _08783_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1036 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15149_ _07795_ _07796_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[7\]
+ VGND VGND VPWR VPWR _07798_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19957_ _01758_ _01755_ _01775_ _10957_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18908_ _11330_ _11331_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[7\]
+ _07816_ VGND VGND VPWR VPWR _11332_ sky130_fd_sc_hd__a2bb2o_1
X_19888_ _01652_ _01673_ _01694_ _01710_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_138_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_218_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18839_ _11232_ _11235_ _11234_ VGND VGND VPWR VPWR _11264_ sky130_fd_sc_hd__o21a_1
XFILLER_0_223_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21850_ _03070_ _03569_ _03570_ _02909_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20801_ _02465_ _02574_ _02575_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21781_ _03503_ _03504_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23520_ clknet_leaf_138_clk _00053_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20732_ _02508_ _02509_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23451_ net392 _04864_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__or2_1
XFILLER_0_212_1097 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20663_ _02436_ _02442_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22402_ _04053_ _04086_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_190_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23382_ net54 _04805_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20594_ _02323_ _02336_ _02375_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22333_ _04017_ _04018_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_1250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22264_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[5\] top_inst.grid_inst.data_path_wires\[18\]\[4\]
+ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24003_ clknet_leaf_82_clk _00536_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[4\]
+ sky130_fd_sc_hd__dfxtp_4
X_21215_ _02927_ _02934_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22195_ _03311_ _03884_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21146_ _02893_ _02021_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__or2_1
XFILLER_0_228_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21077_ _02835_ _02834_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__or2b_1
X_20028_ _01828_ _01830_ _01843_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__a21o_1
XFILLER_0_226_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12850_ _05655_ _05656_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__or2b_1
XFILLER_0_197_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11801_ top_inst.axis_out_inst.out_buff_data\[79\] _04890_ VGND VGND VPWR VPWR _04901_
+ sky130_fd_sc_hd__or2_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _05547_ _05589_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__xnor2_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21979_ top_inst.grid_inst.data_path_wires\[18\]\[4\] VGND VGND VPWR VPWR _03688_
+ sky130_fd_sc_hd__buf_2
XFILLER_0_189_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _07178_ _07211_ _07212_ VGND VGND VPWR VPWR _07213_ sky130_fd_sc_hd__and3_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23718_ clknet_leaf_120_clk _00251_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14451_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[3\]
+ _07060_ _07064_ VGND VGND VPWR VPWR _07146_ sky130_fd_sc_hd__nand4_4
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23649_ clknet_leaf_128_clk net324 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13402_ _06100_ _06154_ _06152_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17170_ _09663_ _09718_ VGND VGND VPWR VPWR _09719_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14382_ _07083_ _07075_ VGND VGND VPWR VPWR _07084_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16121_ net1064 _08183_ _08709_ _08692_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__o211a_1
X_13333_ _06106_ _06107_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1069 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_130_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_130_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_40_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16052_ _08642_ _08644_ _08645_ _08658_ VGND VGND VPWR VPWR _08659_ sky130_fd_sc_hd__o31a_1
XFILLER_0_228_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13264_ _05886_ _06040_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_971 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15003_ _07610_ _07608_ _07629_ _07627_ VGND VGND VPWR VPWR _07657_ sky130_fd_sc_hd__nand4_1
X_12215_ _05044_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__clkbuf_4
X_13195_ _05746_ _05768_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19811_ _01632_ _01636_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_236_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12146_ net463 _05089_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_236_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19742_ _01534_ _01536_ _01535_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_159_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16954_ _09465_ _09508_ VGND VGND VPWR VPWR _09509_ sky130_fd_sc_hd__xor2_2
X_12077_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[5\] _05050_
+ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__or2_1
XFILLER_0_202_1299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15905_ _08490_ _08489_ VGND VGND VPWR VPWR _08516_ sky130_fd_sc_hd__or2b_1
XFILLER_0_217_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19673_ _01500_ net250 _01483_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_205_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16885_ _09439_ _09440_ _09422_ VGND VGND VPWR VPWR _09442_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_1126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18624_ _10840_ _11045_ _11081_ VGND VGND VPWR VPWR _11083_ sky130_fd_sc_hd__nor3_1
XFILLER_0_205_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15836_ _08436_ _08448_ VGND VGND VPWR VPWR _08449_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18555_ _11014_ _11015_ VGND VGND VPWR VPWR _11016_ sky130_fd_sc_hd__and2_1
XFILLER_0_188_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12979_ _05768_ _05294_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__or2_1
XTAP_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ _08369_ _08381_ VGND VGND VPWR VPWR _08382_ sky130_fd_sc_hd__xnor2_1
XTAP_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17506_ _10032_ _10033_ _10034_ _10024_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14718_ _07328_ _07376_ _07375_ VGND VGND VPWR VPWR _07406_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18486_ _10922_ _10948_ VGND VGND VPWR VPWR _10949_ sky130_fd_sc_hd__xor2_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15698_ top_inst.grid_inst.data_path_wires\[7\]\[2\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[5\]
+ VGND VGND VPWR VPWR _08314_ sky130_fd_sc_hd__nand2_1
X_17437_ _09915_ _09973_ VGND VGND VPWR VPWR _09974_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14649_ _07291_ _07294_ VGND VGND VPWR VPWR _07339_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_16 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_27 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17368_ _09880_ _09904_ VGND VGND VPWR VPWR _09908_ sky130_fd_sc_hd__or2b_1
XANTENNA_49 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19107_ _11524_ _11525_ VGND VGND VPWR VPWR _11526_ sky130_fd_sc_hd__nor2_1
X_16319_ _08899_ _08900_ VGND VGND VPWR VPWR _08901_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_121_clk clknet_4_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17299_ _09812_ _09817_ _09840_ _09795_ VGND VGND VPWR VPWR _09843_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19038_ _11457_ _11458_ VGND VGND VPWR VPWR _11459_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput101 net101 VGND VGND VPWR VPWR output_tdata[41] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_242_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput112 net112 VGND VGND VPWR VPWR output_tdata[51] sky130_fd_sc_hd__clkbuf_4
Xoutput123 net123 VGND VGND VPWR VPWR output_tdata[61] sky130_fd_sc_hd__clkbuf_4
Xoutput134 net134 VGND VGND VPWR VPWR output_tdata[71] sky130_fd_sc_hd__buf_2
XFILLER_0_140_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput145 net145 VGND VGND VPWR VPWR output_tdata[81] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput156 net156 VGND VGND VPWR VPWR output_tdata[91] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21000_ _02463_ _02766_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22951_ net704 _04562_ _04563_ _04564_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21902_ _03612_ _03619_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_190_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22882_ top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[6\] _04517_ VGND
+ VGND VPWR VPWR _04525_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24621_ clknet_leaf_21_clk net582 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[97\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21833_ _03553_ _03533_ _03531_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24552_ clknet_leaf_133_clk _01085_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dfxtp_4
X_21764_ _03487_ _03488_ _05732_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__a21o_1
XFILLER_0_176_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23503_ clknet_leaf_140_clk net685 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[93\]
+ sky130_fd_sc_hd__dfxtp_1
X_20715_ _02492_ _02487_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24483_ clknet_leaf_115_clk _01016_ VGND VGND VPWR VPWR top_inst.valid_pipe\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21695_ _03123_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23434_ net964 _04827_ _04838_ _04831_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20646_ _02408_ _02409_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23365_ net46 _04792_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20577_ _01997_ _02229_ _02357_ _02358_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_112_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22316_ _03977_ _04002_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23296_ net140 _04753_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1042 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22247_ _03889_ _03896_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__or2b_1
X_12000_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[4\] _05010_
+ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__or2_1
XFILLER_0_218_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22178_ top_inst.grid_inst.data_path_wires\[18\]\[0\] _03713_ VGND VGND VPWR VPWR
+ _03868_ sky130_fd_sc_hd__and2b_1
XFILLER_0_218_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21129_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _02882_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_233_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13951_ _06669_ _06670_ VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__nor2_1
XFILLER_0_199_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12902_ _05677_ _05680_ _05705_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__nand3_1
XFILLER_0_92_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16670_ _09194_ _09192_ _09197_ _09189_ VGND VGND VPWR VPWR _09233_ sky130_fd_sc_hd__a22o_1
X_13882_ _06618_ _06620_ VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__or2_1
XFILLER_0_202_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12833_ _05267_ top_inst.skew_buff_inst.row\[0\].output_reg\[6\] VGND VGND VPWR VPWR
+ _05640_ sky130_fd_sc_hd__and2b_1
XFILLER_0_9_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15621_ _08135_ _08167_ VGND VGND VPWR VPWR _08239_ sky130_fd_sc_hd__nand2_1
XFILLER_0_198_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18340_ _10802_ _10805_ VGND VGND VPWR VPWR _10806_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _05571_ _05572_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__xnor2_1
X_15552_ net1075 _06660_ _08174_ _08166_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__o211a_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14503_ _07172_ _07173_ _07194_ _07195_ VGND VGND VPWR VPWR _07196_ sky130_fd_sc_hd__a211o_1
XFILLER_0_132_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15483_ _08101_ _08109_ VGND VGND VPWR VPWR _08123_ sky130_fd_sc_hd__or2_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18271_ _10713_ _10714_ _10737_ _10738_ VGND VGND VPWR VPWR _10739_ sky130_fd_sc_hd__a211oi_2
X_12695_ _05455_ _05458_ _05456_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_167_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17222_ net199 _09768_ VGND VGND VPWR VPWR _09769_ sky130_fd_sc_hd__nor2_1
X_14434_ _07118_ _07111_ _07129_ VGND VGND VPWR VPWR _07130_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_830 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput14 input_tdata[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
XFILLER_0_64_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17153_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[14\] _09459_ _09417_
+ VGND VGND VPWR VPWR _09703_ sky130_fd_sc_hd__a21o_1
X_14365_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _07070_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput25 input_tdata[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_4
XFILLER_0_128_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput36 reset VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_103_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16104_ _08673_ _08681_ _08696_ _08692_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__o211a_1
X_13316_ _06089_ _06090_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17084_ _09361_ _09377_ _09215_ net219 VGND VGND VPWR VPWR _09636_ sky130_fd_sc_hd__or4b_1
Xhold809 top_inst.axis_in_inst.inbuf_bus\[17\] VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__dlygate4sd3_1
X_14296_ _06936_ _07004_ VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_896 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13247_ _05977_ _05980_ _05978_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16035_ _08640_ _08641_ VGND VGND VPWR VPWR _08643_ sky130_fd_sc_hd__and2_1
XFILLER_0_243_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13178_ _05908_ _05902_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12129_ net256 _05084_ _05087_ _05088_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__o211a_1
XFILLER_0_237_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17986_ _10457_ _10472_ _10470_ VGND VGND VPWR VPWR _10489_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19725_ _01519_ _01553_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__or2_1
X_16937_ _09453_ _09492_ VGND VGND VPWR VPWR _09493_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_174_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19656_ _01402_ _01484_ _01485_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__or3_4
X_16868_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[3\]
+ net215 _09209_ VGND VGND VPWR VPWR _09425_ sky130_fd_sc_hd__and4_1
XFILLER_0_215_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18607_ _11030_ _11005_ VGND VGND VPWR VPWR _11067_ sky130_fd_sc_hd__and2b_1
X_15819_ _08391_ _08396_ _08432_ VGND VGND VPWR VPWR _08433_ sky130_fd_sc_hd__a21oi_1
X_19587_ _01415_ _01416_ _01417_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16799_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[6\] _09357_ _08307_
+ VGND VGND VPWR VPWR _09358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18538_ _10960_ _10998_ VGND VGND VPWR VPWR _11000_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18469_ _10892_ _10931_ VGND VGND VPWR VPWR _10932_ sky130_fd_sc_hd__nor2_2
XFILLER_0_185_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20500_ _01995_ _02188_ _02283_ _02186_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21480_ _03212_ _03213_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20431_ _02215_ _02216_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__or2b_1
XFILLER_0_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_910 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23150_ net359 _04671_ _04678_ _04675_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20362_ top_inst.grid_inst.data_path_wires\[16\]\[5\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[1\]
+ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22101_ _03786_ _03792_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23081_ net20 _04628_ _04638_ _04632_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__o211a_1
X_20293_ _02079_ _02080_ _02078_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22032_ _03684_ _03700_ _03682_ _03698_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__nand4_1
XTAP_6319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23983_ clknet_leaf_81_clk _00516_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22934_ net590 _04548_ _04554_ _04551_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22865_ net708 _04504_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24604_ clknet_leaf_21_clk _01137_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dfxtp_1
X_21816_ _03514_ _03517_ _03535_ _03496_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_94_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22796_ _04457_ _04464_ _06178_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24535_ clknet_leaf_131_clk _01068_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_52_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21747_ _03447_ _03450_ _03449_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__o21bai_2
XPHY_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24466_ clknet_leaf_57_clk _00999_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12480_ _05300_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21678_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[17\] _03122_ VGND
+ VGND VPWR VPWR _03406_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23417_ top_inst.axis_out_inst.out_buff_data\[98\] _04596_ VGND VGND VPWR VPWR _04829_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20629_ _02408_ _02409_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__xor2_1
X_24397_ clknet_leaf_38_clk net785 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14150_ _06817_ _06818_ _06814_ VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__or3b_1
XFILLER_0_145_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23348_ _04684_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_1125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13101_ net169 _05880_ _05848_ _05844_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14081_ _06717_ _06754_ _06796_ VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__a21o_1
XFILLER_0_162_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23279_ _04684_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_104_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13032_ _05809_ _05814_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__xor2_1
XFILLER_0_219_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17840_ _10333_ _10334_ _10346_ VGND VGND VPWR VPWR _10347_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_219_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17771_ _10271_ _10273_ _10269_ VGND VGND VPWR VPWR _10279_ sky130_fd_sc_hd__a21o_1
X_14983_ _05772_ VGND VGND VPWR VPWR _07641_ sky130_fd_sc_hd__buf_2
XFILLER_0_234_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19510_ _11722_ _01343_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__and2_1
XFILLER_0_195_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16722_ _09280_ _09281_ _09272_ VGND VGND VPWR VPWR _09283_ sky130_fd_sc_hd__a21o_1
X_13934_ _06640_ _06622_ _06637_ _06618_ VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19441_ _01274_ _01275_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__nor2_1
X_16653_ net219 VGND VGND VPWR VPWR _09219_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13865_ _06578_ _06582_ _06604_ _06404_ VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_187_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15604_ _08201_ _08222_ VGND VGND VPWR VPWR _08223_ sky130_fd_sc_hd__xor2_2
X_12816_ _05582_ _05623_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__or2_1
X_19372_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[3\] _01187_ _01188_
+ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_70_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_922 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16584_ _09150_ _09158_ VGND VGND VPWR VPWR _09159_ sky130_fd_sc_hd__xnor2_1
X_13796_ _06458_ net181 _06538_ VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_202_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18323_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[7\] _10755_ _10756_
+ VGND VGND VPWR VPWR _10789_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_151_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15535_ _08143_ _07639_ _08162_ _08142_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12747_ _05554_ _05555_ _05516_ _05518_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__a211o_1
XFILLER_0_167_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18254_ _10717_ _10721_ VGND VGND VPWR VPWR _10722_ sky130_fd_sc_hd__xor2_1
X_12678_ _05304_ _05488_ _05283_ _05302_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__a22o_1
X_15466_ _08102_ _08106_ VGND VGND VPWR VPWR _08107_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17205_ _09417_ _09418_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[17\]
+ VGND VGND VPWR VPWR _09753_ sky130_fd_sc_hd__or3b_1
XFILLER_0_170_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14417_ net173 _07112_ _05315_ VGND VGND VPWR VPWR _07114_ sky130_fd_sc_hd__o21a_1
XFILLER_0_181_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18185_ _10643_ _10635_ _10655_ VGND VGND VPWR VPWR _10656_ sky130_fd_sc_hd__a21o_1
XFILLER_0_231_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15397_ _08038_ _08039_ VGND VGND VPWR VPWR _08040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17136_ _09685_ _09683_ VGND VGND VPWR VPWR _09687_ sky130_fd_sc_hd__or2b_1
XFILLER_0_167_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14348_ _07050_ _07055_ VGND VGND VPWR VPWR _07056_ sky130_fd_sc_hd__nor2_1
Xhold606 top_inst.axis_out_inst.out_buff_data\[116\] VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold617 top_inst.axis_out_inst.out_buff_data\[21\] VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold628 top_inst.axis_out_inst.out_buff_data\[115\] VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14279_ _06956_ VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__inv_2
X_17067_ net1091 _09494_ VGND VGND VPWR VPWR _09620_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_1404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold639 top_inst.axis_out_inst.out_buff_data\[57\] VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16018_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[15\] _07576_ VGND
+ VGND VPWR VPWR _08626_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17969_ _10457_ _10472_ VGND VGND VPWR VPWR _10473_ sky130_fd_sc_hd__xor2_2
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_236_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19708_ _01534_ _01535_ _01536_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__nand3_1
XFILLER_0_100_1178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20980_ _02463_ _02747_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_174_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_1377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19639_ _01467_ _01469_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22650_ _04296_ _04299_ _04321_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_177_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21601_ _03320_ _03331_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__xnor2_2
X_22581_ _04259_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24320_ clknet_leaf_143_clk _00853_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[95\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21532_ _03251_ _03264_ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__xor2_1
XFILLER_0_173_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24251_ clknet_leaf_107_clk _00784_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21463_ _03154_ _03189_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23202_ net95 _04701_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__or2_1
XFILLER_0_181_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20414_ _02197_ _02198_ _02191_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__a21o_1
X_24182_ clknet_leaf_29_clk _00715_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[25\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21394_ _03124_ _03129_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23133_ net755 _04656_ _04668_ _04662_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20345_ _02099_ _02131_ _05335_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23064_ _04602_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__buf_2
XFILLER_0_102_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20276_ _02063_ _02064_ _02065_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__and3_2
XFILLER_0_12_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22015_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _03713_ sky130_fd_sc_hd__clkbuf_4
XTAP_6149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ top_inst.axis_out_inst.out_buff_data\[60\] _04996_ VGND VGND VPWR VPWR _05003_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_242_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23966_ clknet_leaf_85_clk _00499_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_231_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22917_ net389 _04535_ _04544_ _04537_ VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__o211a_1
X_23897_ clknet_leaf_52_clk _00430_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22848_ net850 _04496_ _04505_ _04498_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13650_ _06347_ _06341_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__or2b_1
XFILLER_0_196_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ _05302_ _05298_ _05272_ _05279_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__nand4_2
X_13581_ top_inst.grid_inst.data_path_wires\[2\]\[0\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__or2b_1
XFILLER_0_13_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22779_ _04446_ _04447_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12532_ _05283_ _05322_ _05334_ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__o21bai_1
X_15320_ _07956_ _07964_ VGND VGND VPWR VPWR _07965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_1203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24518_ clknet_leaf_135_clk _01051_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dfxtp_2
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12463_ _05286_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__buf_2
XFILLER_0_164_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15251_ _07896_ _07897_ VGND VGND VPWR VPWR _07898_ sky130_fd_sc_hd__xnor2_1
X_24449_ clknet_leaf_63_clk _00982_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_14202_ _06872_ _06874_ VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15182_ _07781_ _07782_ _07829_ VGND VGND VPWR VPWR _07830_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_22_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12394_ net567 _05230_ _05239_ _05234_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14133_ _05632_ _06847_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19990_ _01806_ _01807_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__xor2_1
XFILLER_0_205_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14064_ _06778_ _06779_ VGND VGND VPWR VPWR _06780_ sky130_fd_sc_hd__nand2_1
X_18941_ _11307_ _11321_ _11363_ VGND VGND VPWR VPWR _11364_ sky130_fd_sc_hd__o21a_1
XFILLER_0_162_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13015_ _05785_ _05797_ _05798_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__nor3_1
XFILLER_0_24_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18872_ _11296_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_1410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17823_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[10\] _10236_ VGND
+ VGND VPWR VPWR _10330_ sky130_fd_sc_hd__xnor2_2
XTAP_6683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17754_ _10218_ _10195_ VGND VGND VPWR VPWR _10263_ sky130_fd_sc_hd__or2b_1
XFILLER_0_221_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14966_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _07629_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1040 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16705_ _05787_ VGND VGND VPWR VPWR _09266_ sky130_fd_sc_hd__buf_6
X_13917_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _06645_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_221_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17685_ _10167_ _10176_ _10178_ VGND VGND VPWR VPWR _10195_ sky130_fd_sc_hd__o21ai_1
X_14897_ _07561_ _07563_ VGND VGND VPWR VPWR _07580_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19424_ _01250_ _01251_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__nand2_1
X_16636_ top_inst.skew_buff_inst.row\[2\].output_reg\[4\] top_inst.axis_in_inst.inbuf_bus\[20\]
+ _05265_ VGND VGND VPWR VPWR _09205_ sky130_fd_sc_hd__mux2_4
XFILLER_0_212_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13848_ _06527_ _06558_ _06559_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_57_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19355_ _01191_ _01192_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__or2b_1
XFILLER_0_9_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16567_ _09141_ _09142_ VGND VGND VPWR VPWR _09143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13779_ _06515_ _06517_ VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__or2_1
XFILLER_0_169_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18306_ _10766_ _10772_ VGND VGND VPWR VPWR _10773_ sky130_fd_sc_hd__xor2_2
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15518_ _08150_ _08140_ VGND VGND VPWR VPWR _08151_ sky130_fd_sc_hd__or2_1
X_19286_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _11688_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16498_ _09072_ _09074_ _05353_ VGND VGND VPWR VPWR _09076_ sky130_fd_sc_hd__a21o_1
X_18237_ _10703_ _10705_ VGND VGND VPWR VPWR _10706_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15449_ _08088_ _08090_ VGND VGND VPWR VPWR _08091_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18168_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[2\] _10639_ VGND
+ VGND VPWR VPWR _10640_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold403 top_inst.deskew_buff_inst.col_input\[7\] VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__dlygate4sd3_1
X_17119_ _09667_ _09669_ VGND VGND VPWR VPWR _09670_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold414 top_inst.deskew_buff_inst.col_input\[13\] VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 _00966_ VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18099_ _10585_ _08674_ VGND VGND VPWR VPWR _10586_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold436 top_inst.axis_out_inst.out_buff_data\[12\] VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold447 top_inst.axis_out_inst.out_buff_data\[87\] VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__dlygate4sd3_1
X_20130_ _01918_ _01933_ _01941_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__a21oi_1
Xhold458 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[16\] VGND
+ VGND VPWR VPWR net640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 top_inst.axis_out_inst.out_buff_data\[47\] VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap177 _02279_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__buf_1
XFILLER_0_229_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_1267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20061_ _01871_ _01875_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__xor2_2
XFILLER_0_239_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23820_ clknet_leaf_93_clk _00353_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23751_ clknet_leaf_135_clk net299 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_20963_ _02730_ _02731_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__nand2_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_92_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22702_ _04374_ _04366_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__xnor2_1
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23682_ clknet_leaf_117_clk net312 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20894_ _02653_ _02654_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22633_ _04061_ _04308_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22564_ _04092_ _04241_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24303_ clknet_leaf_2_clk _00836_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[78\]
+ sky130_fd_sc_hd__dfxtp_1
X_21515_ _03246_ _03247_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__xor2_1
X_22495_ _04174_ _04176_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24234_ clknet_leaf_112_clk _00767_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_21446_ _03141_ _03143_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_224_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24165_ clknet_leaf_9_clk _00698_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_102_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21377_ net808 _02638_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23116_ _04658_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__buf_2
X_20328_ _02112_ _02113_ _02114_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__a21o_1
X_24096_ clknet_leaf_99_clk _00629_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_23047_ net965 _04616_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20259_ _02033_ _02046_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__nand2_1
XTAP_5212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14820_ _07493_ _07494_ _07504_ VGND VGND VPWR VPWR _07506_ sky130_fd_sc_hd__nand3_1
XFILLER_0_200_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_203_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ _05633_ VGND VGND VPWR VPWR _07439_ sky130_fd_sc_hd__clkbuf_8
XTAP_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23949_ clknet_leaf_81_clk _00482_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11963_ top_inst.axis_out_inst.out_buff_data\[53\] _04982_ VGND VGND VPWR VPWR _04993_
+ sky130_fd_sc_hd__or2_1
XTAP_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_83_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_16
XTAP_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _06439_ _06441_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__or2_1
X_17470_ _10001_ _09995_ _10004_ VGND VGND VPWR VPWR _10006_ sky130_fd_sc_hd__nand3_1
XFILLER_0_170_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14682_ _07365_ _07370_ VGND VGND VPWR VPWR _07371_ sky130_fd_sc_hd__xor2_1
XTAP_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11894_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[23\] _04943_
+ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16421_ _08986_ _08988_ VGND VGND VPWR VPWR _09000_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13633_ _06374_ _06379_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19140_ top_inst.grid_inst.data_path_wires\[13\]\[7\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _11558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16352_ _08931_ _08932_ VGND VGND VPWR VPWR _08933_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13564_ _06304_ _06312_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__xnor2_2
X_15303_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[11\] VGND VGND
+ VPWR VPWR _07948_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12515_ _05330_ _05331_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__xnor2_1
X_19071_ _11488_ _11490_ VGND VGND VPWR VPWR _11491_ sky130_fd_sc_hd__xor2_1
XFILLER_0_136_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16283_ _08864_ _08865_ VGND VGND VPWR VPWR _08866_ sky130_fd_sc_hd__nor2_1
X_13495_ top_inst.grid_inst.data_path_wires\[2\]\[3\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[2\]\[4\]
+ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18022_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[15\] _10367_ VGND
+ VGND VPWR VPWR _10524_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12446_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _05273_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_151_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15234_ top_inst.grid_inst.data_path_wires\[6\]\[7\] _07631_ VGND VGND VPWR VPWR
+ _07881_ sky130_fd_sc_hd__nand2_4
XFILLER_0_129_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1088 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15165_ _07812_ _07813_ VGND VGND VPWR VPWR _07814_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12377_ net896 _05217_ _05229_ _05221_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__o211a_1
XFILLER_0_244_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14116_ _06827_ _06828_ _06830_ VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__a21boi_1
X_19973_ _01790_ _01791_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__nor2_1
X_15096_ _07608_ top_inst.grid_inst.data_path_wires\[6\]\[0\] _07640_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[5\]
+ VGND VGND VPWR VPWR _07746_ sky130_fd_sc_hd__nand4_2
XFILLER_0_120_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18924_ _11145_ _11154_ _11344_ _11345_ VGND VGND VPWR VPWR _11347_ sky130_fd_sc_hd__nand4_1
X_14047_ _06704_ _06728_ _06727_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_226_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18855_ _11274_ _11279_ VGND VGND VPWR VPWR _11280_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_235_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17806_ _10282_ _10313_ VGND VGND VPWR VPWR _10314_ sky130_fd_sc_hd__xor2_1
XFILLER_0_237_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18786_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[4\] _11212_ VGND
+ VGND VPWR VPWR _11213_ sky130_fd_sc_hd__xor2_4
XFILLER_0_59_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15998_ _08605_ _08606_ VGND VGND VPWR VPWR _08607_ sky130_fd_sc_hd__nor2_1
XFILLER_0_222_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_221_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17737_ top_inst.grid_inst.data_path_wires\[11\]\[1\] VGND VGND VPWR VPWR _10246_
+ sky130_fd_sc_hd__inv_2
X_14949_ _04868_ VGND VGND VPWR VPWR _07617_ sky130_fd_sc_hd__buf_4
XFILLER_0_222_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_74_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_106_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17668_ _10166_ _10177_ VGND VGND VPWR VPWR _10179_ sky130_fd_sc_hd__or2_1
XFILLER_0_202_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19407_ _11701_ _11677_ _01240_ _01241_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_106_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16619_ top_inst.skew_buff_inst.row\[2\].output_reg\[1\] top_inst.axis_in_inst.inbuf_bus\[17\]
+ _07059_ VGND VGND VPWR VPWR _09191_ sky130_fd_sc_hd__mux2_4
XFILLER_0_119_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17599_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[3\] _10091_ _10092_
+ VGND VGND VPWR VPWR _10112_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19338_ _11724_ _11731_ VGND VGND VPWR VPWR _11732_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19269_ net1057 _11662_ _11675_ VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21300_ _02875_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[1\] _02882_
+ _02878_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22280_ _03936_ _03967_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold200 top_inst.axis_out_inst.out_buff_data\[20\] VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__dlygate4sd3_1
X_21231_ _02965_ _02970_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__xnor2_2
Xhold211 top_inst.axis_out_inst.out_buff_data\[84\] VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold222 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[7\] VGND VGND
+ VPWR VPWR net404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 top_inst.axis_out_inst.out_buff_data\[89\] VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 top_inst.deskew_buff_inst.col_input\[10\] VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 top_inst.deskew_buff_inst.col_input\[15\] VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__dlygate4sd3_1
X_21162_ _02904_ _02905_ _02899_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold266 _00136_ VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold277 _00141_ VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__dlygate4sd3_1
X_20113_ _01924_ _01925_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__and2_1
Xhold288 _00156_ VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[2\] VGND
+ VGND VPWR VPWR net481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21093_ _02460_ _02841_ _02528_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20044_ _01834_ _01859_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_176_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23803_ clknet_leaf_77_clk _00336_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ _03680_ _02881_ _03699_ _03660_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_65_clk clknet_4_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 _05275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_241_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_117 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20946_ _02710_ _02712_ _02714_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__nor3_1
X_23734_ clknet_leaf_125_clk _00267_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23665_ clknet_leaf_132_clk net384 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20877_ _02617_ _02648_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22616_ _04288_ _04292_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__xor2_2
XFILLER_0_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23596_ clknet_leaf_100_clk _00129_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22547_ _04225_ _04226_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12300_ net600 _05178_ _05186_ _05182_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13280_ _06050_ _06054_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22478_ _04118_ _04151_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12231_ net528 _05143_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__or2_1
XFILLER_0_228_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24217_ clknet_leaf_118_clk _00750_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_21429_ _02878_ _02887_ _03131_ _03132_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24148_ clknet_leaf_16_clk _00681_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[13\]\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_47_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12162_ top_inst.axis_out_inst.out_buff_data\[10\] _05102_ VGND VGND VPWR VPWR _05107_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_130_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_562 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16970_ _09481_ _09500_ _09523_ _09524_ VGND VGND VPWR VPWR _09525_ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_1284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12093_ net1106 _05063_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__or2_1
X_24079_ clknet_leaf_113_clk _00612_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15921_ _08409_ _08482_ _08444_ VGND VGND VPWR VPWR _08532_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_198_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_975 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18640_ _10933_ VGND VGND VPWR VPWR _11098_ sky130_fd_sc_hd__inv_2
XTAP_5075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15852_ _08424_ _08425_ _08464_ VGND VGND VPWR VPWR _08465_ sky130_fd_sc_hd__o21a_1
XFILLER_0_232_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _07450_ _07488_ VGND VGND VPWR VPWR _07489_ sky130_fd_sc_hd__nor2_1
XFILLER_0_203_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ _10964_ _10993_ _10991_ VGND VGND VPWR VPWR _11032_ sky130_fd_sc_hd__o21a_1
XTAP_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15783_ _08387_ _08389_ VGND VGND VPWR VPWR _08397_ sky130_fd_sc_hd__or2_1
XFILLER_0_235_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_157_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12995_ net1060 _05314_ _05780_ _05767_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__o211a_1
XTAP_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17522_ _10025_ _08681_ _10045_ _10024_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__o211a_1
XTAP_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14734_ _07379_ _07381_ VGND VGND VPWR VPWR _07422_ sky130_fd_sc_hd__nand2_1
XTAP_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ top_inst.axis_out_inst.out_buff_data\[45\] _04982_ VGND VGND VPWR VPWR _04984_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ _09892_ _09987_ _09989_ VGND VGND VPWR VPWR _09990_ sky130_fd_sc_hd__a21oi_2
X_14665_ _07316_ _07354_ VGND VGND VPWR VPWR _07355_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[15\] _04943_
+ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__or2_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16404_ _08981_ _08983_ VGND VGND VPWR VPWR _08984_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13616_ _06363_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__clkbuf_1
X_17384_ _09877_ _09920_ _09923_ VGND VGND VPWR VPWR _09924_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14596_ _07079_ _07074_ _07078_ _07082_ VGND VGND VPWR VPWR _07287_ sky130_fd_sc_hd__and4_1
XFILLER_0_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19123_ _11540_ _11541_ VGND VGND VPWR VPWR _11542_ sky130_fd_sc_hd__nor2_1
X_16335_ _08872_ _08916_ VGND VGND VPWR VPWR _08917_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13547_ _06184_ top_inst.grid_inst.data_path_wires\[2\]\[0\] _06214_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[5\]
+ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__nand4_2
XFILLER_0_171_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19054_ _11472_ _11471_ VGND VGND VPWR VPWR _11474_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16266_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[7\] _08847_ _08848_
+ VGND VGND VPWR VPWR _08849_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13478_ top_inst.grid_inst.data_path_wires\[2\]\[1\] top_inst.grid_inst.data_path_wires\[2\]\[0\]
+ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[3\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[2\]
+ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__and4_1
XFILLER_0_242_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18005_ _10489_ _10507_ VGND VGND VPWR VPWR _10508_ sky130_fd_sc_hd__or2b_1
XFILLER_0_129_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15217_ _07820_ _07864_ VGND VGND VPWR VPWR _07865_ sky130_fd_sc_hd__xor2_1
X_12429_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[29\] _05248_
+ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16197_ _08747_ _08748_ _08781_ VGND VGND VPWR VPWR _08782_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15148_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[7\] _07795_ _07796_
+ VGND VGND VPWR VPWR _07797_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19956_ _01758_ _01755_ _01775_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__a21oi_1
X_15079_ _07671_ _07692_ VGND VGND VPWR VPWR _07730_ sky130_fd_sc_hd__nor2_1
XFILLER_0_177_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18907_ _11328_ _11329_ _05353_ VGND VGND VPWR VPWR _11331_ sky130_fd_sc_hd__a21o_1
X_19887_ _01678_ _01671_ _01693_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_207_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_0__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_4_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_18838_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[5\] _11240_ _11241_
+ VGND VGND VPWR VPWR _11263_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_101_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18769_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[3\] _11195_ _11196_
+ VGND VGND VPWR VPWR _11197_ sky130_fd_sc_hd__and3_1
XFILLER_0_179_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_47_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_223_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20800_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[18\] _02467_ VGND
+ VGND VPWR VPWR _02575_ sky130_fd_sc_hd__or2_1
XFILLER_0_222_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21780_ _03501_ _03502_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__and2_1
XFILLER_0_194_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1010 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20731_ _02506_ _02507_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__and2_1
XFILLER_0_175_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23450_ net508 _04840_ _04847_ _04844_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20662_ _02437_ _02441_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22401_ _04054_ _04085_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23381_ net392 _04804_ _04810_ _04808_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20593_ _02334_ _02335_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22332_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[11\] _03893_ VGND
+ VGND VPWR VPWR _04018_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_190_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22263_ _03949_ _03950_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24002_ clknet_leaf_46_clk _00535_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_21214_ _02950_ _02954_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__xor2_2
X_22194_ _03882_ _03883_ top_inst.deskew_buff_inst.col_input\[103\] _05354_ VGND VGND
+ VPWR VPWR _03884_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_112_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21145_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _02893_ sky130_fd_sc_hd__buf_2
XFILLER_0_217_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_217_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21076_ net327 _02491_ _02838_ _02839_ _01863_ VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__o221a_1
XFILLER_0_233_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20027_ _01563_ _01829_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_241_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_38_clk clknet_4_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11800_ net570 _04898_ _04900_ _04889_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__o211a_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12780_ _05587_ _05588_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21978_ _02868_ _02877_ _03687_ _03660_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__o211a_1
Xrebuffer70 _09560_ VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23717_ clknet_leaf_121_clk _00250_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20929_ _02667_ _02697_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__nand2_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14450_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[2\] _07069_ VGND
+ VGND VPWR VPWR _07145_ sky130_fd_sc_hd__nand2_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23648_ clknet_leaf_127_clk _00181_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13401_ _06113_ _06158_ _06156_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__a21oi_1
X_14381_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _07083_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23579_ clknet_leaf_106_clk _00112_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16120_ _08707_ _08708_ _06682_ VGND VGND VPWR VPWR _08709_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13332_ _06104_ _06105_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16051_ _08642_ _08657_ VGND VGND VPWR VPWR _08658_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13263_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[10\] _05354_ _06038_
+ _06039_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_983 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15002_ _07608_ _07629_ _07627_ _07610_ VGND VGND VPWR VPWR _07656_ sky130_fd_sc_hd__a22o_1
X_12214_ net917 _05123_ _05136_ _05128_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__o211a_1
X_13194_ _05970_ _05971_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__nor2_1
XFILLER_0_209_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19810_ _01633_ _01635_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__xnor2_1
X_12145_ _05044_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_236_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16953_ _09207_ _09506_ _09507_ VGND VGND VPWR VPWR _09508_ sky130_fd_sc_hd__a21bo_1
X_19741_ _01566_ _01568_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__xor2_2
X_12076_ _05044_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__buf_2
XFILLER_0_236_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15904_ _05632_ _08515_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__nor2_1
X_19672_ _01483_ _01500_ _01501_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__and3_1
X_16884_ _09422_ _09439_ _09440_ VGND VGND VPWR VPWR _09441_ sky130_fd_sc_hd__and3_1
XFILLER_0_159_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18623_ _10840_ _11045_ _11081_ VGND VGND VPWR VPWR _11082_ sky130_fd_sc_hd__o21a_1
XFILLER_0_235_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_635 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15835_ _08443_ _08447_ VGND VGND VPWR VPWR _08448_ sky130_fd_sc_hd__xor2_1
XFILLER_0_91_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_clk clknet_4_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_16
XTAP_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18554_ _10591_ _10857_ _11013_ VGND VGND VPWR VPWR _11015_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_220_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15766_ _08379_ _08380_ VGND VGND VPWR VPWR _08381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12978_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _05768_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17505_ _10030_ _09206_ VGND VGND VPWR VPWR _10034_ sky130_fd_sc_hd__or2_1
XTAP_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14717_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[10\] _07364_ _07280_
+ VGND VGND VPWR VPWR _07405_ sky130_fd_sc_hd__a21o_1
X_11929_ net845 _04969_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__or2_1
X_18485_ _10946_ _10947_ VGND VGND VPWR VPWR _10948_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15697_ _08311_ _08312_ VGND VGND VPWR VPWR _08313_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17436_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[27\] _09628_ _09629_
+ VGND VGND VPWR VPWR _09973_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14648_ _07336_ _07337_ VGND VGND VPWR VPWR _07338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_17 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_28 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17367_ _08870_ _09906_ _09907_ _09231_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_39 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14579_ _07117_ _07270_ VGND VGND VPWR VPWR _07271_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19106_ _11522_ _11523_ _11520_ VGND VGND VPWR VPWR _11525_ sky130_fd_sc_hd__o21a_1
X_16318_ _08840_ _08842_ _08898_ VGND VGND VPWR VPWR _08900_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17298_ _09833_ _09841_ VGND VGND VPWR VPWR _09842_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19037_ _11428_ _11429_ _11456_ VGND VGND VPWR VPWR _11458_ sky130_fd_sc_hd__nand3_1
XFILLER_0_24_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16249_ _08799_ _08804_ VGND VGND VPWR VPWR _08832_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput102 net102 VGND VGND VPWR VPWR output_tdata[42] sky130_fd_sc_hd__clkbuf_4
Xoutput113 net113 VGND VGND VPWR VPWR output_tdata[52] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_203_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput124 net124 VGND VGND VPWR VPWR output_tdata[62] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput135 net135 VGND VGND VPWR VPWR output_tdata[72] sky130_fd_sc_hd__buf_2
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput146 net146 VGND VGND VPWR VPWR output_tdata[82] sky130_fd_sc_hd__clkbuf_4
Xoutput157 net157 VGND VGND VPWR VPWR output_tdata[92] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_227_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19939_ _01746_ _01747_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__or2b_1
X_22950_ _04550_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21901_ _03618_ _03617_ _03598_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22881_ net828 _04522_ _04523_ _04524_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24620_ clknet_leaf_32_clk _01153_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[96\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21832_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[21\] _03421_ _03422_
+ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24551_ clknet_leaf_103_clk _01084_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dfxtp_2
X_21763_ _03469_ _03486_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23502_ clknet_leaf_141_clk _00035_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[92\]
+ sky130_fd_sc_hd__dfxtp_1
X_20714_ _02457_ _02485_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24482_ clknet_leaf_115_clk _01015_ VGND VGND VPWR VPWR top_inst.valid_pipe\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_21694_ _03376_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__buf_4
XFILLER_0_18_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23433_ net697 _04835_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20645_ _02395_ _02402_ _02424_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23364_ net443 _04791_ _04800_ _04795_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__o211a_1
X_20576_ _02004_ _02015_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[11\]
+ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__and3_1
XFILLER_0_225_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22315_ _03999_ _04001_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__xor2_2
XFILLER_0_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23295_ net705 _04752_ _04761_ _04756_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__o211a_1
XFILLER_0_225_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22246_ _03918_ _03888_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__or2b_1
XFILLER_0_42_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1054 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22177_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[6\] top_inst.grid_inst.data_path_wires\[18\]\[1\]
+ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_178_1008 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21128_ _05269_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_1311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13950_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[3\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[2\]
+ _06622_ top_inst.grid_inst.data_path_wires\[3\]\[0\] VGND VGND VPWR VPWR _06670_
+ sky130_fd_sc_hd__and4_1
X_21059_ _02810_ _02823_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12901_ _05677_ _05680_ _05705_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13881_ _06619_ VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__buf_2
XFILLER_0_9_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15620_ _08225_ _08229_ VGND VGND VPWR VPWR _08238_ sky130_fd_sc_hd__and2b_1
XFILLER_0_236_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12832_ _05304_ _05597_ _05301_ _05302_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _08172_ _08173_ _05336_ VGND VGND VPWR VPWR _08174_ sky130_fd_sc_hd__o21ai_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _05530_ _05531_ _05529_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__o21a_1
XFILLER_0_189_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14502_ _07192_ _07193_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[6\]
+ VGND VGND VPWR VPWR _07195_ sky130_fd_sc_hd__a21oi_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18270_ _10735_ _10736_ _10715_ VGND VGND VPWR VPWR _10738_ sky130_fd_sc_hd__a21oi_1
X_15482_ _08100_ _08122_ _04870_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__o21a_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _05502_ _05504_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__xor2_2
XFILLER_0_182_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17221_ _09743_ _09764_ VGND VGND VPWR VPWR _09768_ sky130_fd_sc_hd__or2b_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14433_ _07125_ _07128_ VGND VGND VPWR VPWR _07129_ sky130_fd_sc_hd__xor2_1
XFILLER_0_193_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17152_ _09678_ _09677_ VGND VGND VPWR VPWR _09702_ sky130_fd_sc_hd__nor2_1
X_14364_ _07068_ VGND VGND VPWR VPWR _07069_ sky130_fd_sc_hd__buf_6
XFILLER_0_182_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput15 input_tdata[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput26 input_tdata[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_123_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16103_ _08695_ _08684_ VGND VGND VPWR VPWR _08696_ sky130_fd_sc_hd__or2_1
X_13315_ _06044_ _06047_ _06045_ VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__o21ba_1
X_17083_ _09597_ _09599_ _09598_ VGND VGND VPWR VPWR _09635_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14295_ _06936_ _07004_ VGND VGND VPWR VPWR _07005_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_1192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16034_ _08614_ _08616_ _08640_ _08641_ VGND VGND VPWR VPWR _08642_ sky130_fd_sc_hd__and4bb_1
X_13246_ _06021_ _06022_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_1034 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_209_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13177_ _05953_ _05955_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12128_ _04994_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__clkbuf_4
X_17985_ _10487_ VGND VGND VPWR VPWR _10488_ sky130_fd_sc_hd__inv_2
XFILLER_0_229_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16936_ _09454_ _09491_ VGND VGND VPWR VPWR _09492_ sky130_fd_sc_hd__xnor2_2
X_19724_ _01520_ _01552_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__xor2_1
X_12059_ _04994_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__buf_2
XFILLER_0_205_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16867_ _09207_ _09206_ _09210_ _09203_ VGND VGND VPWR VPWR _09424_ sky130_fd_sc_hd__a22oi_1
X_19655_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[3\]
+ _11709_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_220_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18606_ _11029_ VGND VGND VPWR VPWR _11066_ sky130_fd_sc_hd__inv_2
X_15818_ _08397_ _08431_ VGND VGND VPWR VPWR _08432_ sky130_fd_sc_hd__xor2_2
XFILLER_0_172_1152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19586_ _01415_ net1126 _01417_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__nand3_4
X_16798_ _09354_ _09356_ VGND VGND VPWR VPWR _09357_ sky130_fd_sc_hd__xor2_1
XFILLER_0_189_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18537_ _10960_ _10998_ VGND VGND VPWR VPWR _10999_ sky130_fd_sc_hd__nand2_1
X_15749_ _08150_ _08159_ _08361_ _08362_ VGND VGND VPWR VPWR _08364_ sky130_fd_sc_hd__nand4_4
XFILLER_0_181_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18468_ _10608_ _10604_ _10595_ VGND VGND VPWR VPWR _10931_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_111_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17419_ _09936_ _09956_ VGND VGND VPWR VPWR _09957_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_173_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18399_ _10847_ _10848_ _10863_ VGND VGND VPWR VPWR _10864_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20430_ _02212_ _02213_ _02214_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__or3b_1
XFILLER_0_172_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20361_ _02144_ _02147_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_9_clk clknet_4_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22100_ _03787_ _03791_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23080_ net1114 _04629_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__or2_1
XFILLER_0_222_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20292_ _02078_ _02079_ _02080_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__nand3_1
XFILLER_0_141_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22031_ _03700_ _03682_ _03698_ _03684_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__a22o_1
XTAP_6309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23982_ clknet_leaf_87_clk _00515_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_138_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22933_ top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[4\] _04543_ VGND
+ VGND VPWR VPWR _04554_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22864_ net1003 _04509_ _04514_ _04511_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24603_ clknet_leaf_30_clk _01136_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_210_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21815_ _03529_ _03536_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__xor2_1
XFILLER_0_167_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22795_ _04364_ _04459_ _04461_ _04463_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__a211o_1
XFILLER_0_151_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24534_ clknet_leaf_131_clk _01067_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dfxtp_2
XPHY_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21746_ _03428_ _03470_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_241_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24465_ clknet_leaf_57_clk _00998_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21677_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[16\] _03376_ _03123_
+ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_93_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23416_ net581 _04827_ _04828_ _04819_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20628_ _02365_ _02370_ _02364_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__a21o_1
X_24396_ clknet_leaf_38_clk net297 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23347_ net993 _04778_ _04790_ _04782_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__o211a_1
X_20559_ _02312_ _02341_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13100_ _05848_ _05844_ net169 _05880_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_46_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14080_ _06750_ _06753_ VGND VGND VPWR VPWR _06796_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23278_ net690 _04739_ _04751_ _04743_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__o211a_1
X_13031_ _05810_ _05813_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__xor2_1
X_22229_ _03915_ _03917_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_203_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17770_ _10262_ _10265_ VGND VGND VPWR VPWR _10278_ sky130_fd_sc_hd__nor2_1
X_14982_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _07640_ sky130_fd_sc_hd__buf_2
XFILLER_0_121_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_238_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16721_ _09272_ _09280_ _09281_ VGND VGND VPWR VPWR _09282_ sky130_fd_sc_hd__nand3_4
X_13933_ net1078 _05788_ _06655_ _06639_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19440_ _11703_ _11701_ net243 _11682_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_1135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16652_ _09217_ VGND VGND VPWR VPWR _09218_ sky130_fd_sc_hd__buf_6
XFILLER_0_134_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13864_ _06578_ _06582_ _06604_ VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15603_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[4\] _08221_ VGND
+ VGND VPWR VPWR _08222_ sky130_fd_sc_hd__xor2_2
XFILLER_0_215_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12815_ _05621_ _05622_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__xor2_1
X_19371_ _01205_ _01206_ _01185_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_187_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16583_ _09156_ _09157_ VGND VGND VPWR VPWR _09158_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13795_ _06202_ _06200_ _06198_ VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18322_ _10753_ _10759_ _10787_ VGND VGND VPWR VPWR _10788_ sky130_fd_sc_hd__a21o_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ _08161_ _07641_ VGND VGND VPWR VPWR _08162_ sky130_fd_sc_hd__or2_1
X_12746_ _05516_ _05518_ _05554_ _05555_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_84_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[6\] _10720_ VGND
+ VGND VPWR VPWR _10721_ sky130_fd_sc_hd__xor2_1
XFILLER_0_194_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15465_ _08103_ _08105_ VGND VGND VPWR VPWR _08106_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12677_ _05278_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17204_ _09588_ _09729_ VGND VGND VPWR VPWR _09752_ sky130_fd_sc_hd__and2_1
X_14416_ net173 _07112_ VGND VGND VPWR VPWR _07113_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18184_ _10647_ _10654_ VGND VGND VPWR VPWR _10655_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15396_ _07956_ _08037_ VGND VGND VPWR VPWR _08039_ sky130_fd_sc_hd__or2_1
X_17135_ _09683_ _09685_ VGND VGND VPWR VPWR _09686_ sky130_fd_sc_hd__or2b_1
XFILLER_0_163_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14347_ _07051_ _07054_ VGND VGND VPWR VPWR _07055_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_170_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold607 top_inst.axis_out_inst.out_buff_data\[34\] VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold618 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[19\] VGND
+ VGND VPWR VPWR net800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17066_ _09583_ _09618_ VGND VGND VPWR VPWR _09619_ sky130_fd_sc_hd__xor2_1
Xhold629 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[18\] VGND
+ VGND VPWR VPWR net811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14278_ _06987_ _06988_ VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16017_ _08625_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__clkbuf_1
X_13229_ _05975_ _05974_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__or2b_1
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17968_ _10470_ _10471_ VGND VGND VPWR VPWR _10472_ sky130_fd_sc_hd__nand2_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19707_ _01298_ _11700_ _11705_ _11703_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_139_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16919_ _09428_ _09430_ _09429_ VGND VGND VPWR VPWR _09475_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17899_ _10324_ _10359_ _10400_ _10403_ _10399_ VGND VGND VPWR VPWR _10404_ sky130_fd_sc_hd__a32o_1
XFILLER_0_205_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19638_ _01345_ _01384_ _01429_ _01468_ _01428_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__o32a_1
XFILLER_0_36_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19569_ _01397_ _01400_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__xor2_1
XFILLER_0_149_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21600_ _03322_ _03330_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__xor2_2
XFILLER_0_192_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22580_ _07707_ _04258_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21531_ _03261_ _03263_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24250_ clknet_leaf_108_clk _00783_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_21462_ _03196_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_173_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23201_ net844 _04700_ _04708_ _04704_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__o211a_1
X_20413_ _02191_ _02197_ _02198_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__nand3_1
XFILLER_0_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24181_ clknet_leaf_29_clk _00714_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_21393_ _03125_ _03128_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23132_ net143 _04659_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__or2_1
X_20344_ _02099_ _02131_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__and2_1
XFILLER_0_226_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23063_ _04600_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20275_ _02007_ _02028_ _02042_ _02044_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__a31o_1
XFILLER_0_222_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22014_ _03693_ _05270_ _03712_ _03702_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__o211a_1
XTAP_6139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23965_ clknet_leaf_89_clk _00498_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_216_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22916_ top_inst.skew_buff_inst.row\[2\].output_reg\[5\] _04543_ VGND VGND VPWR VPWR
+ _04544_ sky130_fd_sc_hd__or2_1
X_23896_ clknet_leaf_52_clk _00429_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22847_ top_inst.skew_buff_inst.row\[3\].output_reg\[7\] _04504_ VGND VGND VPWR VPWR
+ _04505_ sky130_fd_sc_hd__or2_1
XFILLER_0_196_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12600_ _05302_ _05272_ _05279_ _05298_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__a22o_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_233_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13580_ top_inst.grid_inst.data_path_wires\[2\]\[1\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22778_ _04390_ _04445_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12531_ _05345_ _05346_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__and2_1
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24517_ clknet_leaf_135_clk _01050_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_54_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21729_ _03452_ _03454_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__xor2_1
XFILLER_0_192_950 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15250_ _07847_ _07850_ VGND VGND VPWR VPWR _07897_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12462_ top_inst.skew_buff_inst.row\[0\].output_reg\[3\] top_inst.axis_in_inst.inbuf_bus\[3\]
+ net211 VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__mux2_4
X_24448_ clknet_leaf_63_clk net259 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[0\].output_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14201_ _06869_ _06913_ VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15181_ _07783_ _07784_ VGND VGND VPWR VPWR _07829_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24379_ clknet_leaf_37_clk _00912_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12393_ net566 _05235_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14132_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[8\] _05634_ _06845_
+ _06846_ VGND VGND VPWR VPWR _06847_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14063_ _06630_ _06643_ _06776_ _06777_ VGND VGND VPWR VPWR _06779_ sky130_fd_sc_hd__nand4_2
X_18940_ _11308_ _11320_ VGND VGND VPWR VPWR _11363_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13014_ _05741_ _05775_ _05777_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__nor3_1
XFILLER_0_219_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18871_ _10641_ _11295_ VGND VGND VPWR VPWR _11296_ sky130_fd_sc_hd__and2_1
XTAP_6640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17822_ _10040_ _10047_ _10292_ _10293_ VGND VGND VPWR VPWR _10329_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14965_ _07606_ _06647_ _07628_ _07618_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__o211a_1
X_17753_ _10231_ _10261_ VGND VGND VPWR VPWR _10262_ sky130_fd_sc_hd__xnor2_1
XTAP_5994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16704_ _09265_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__clkbuf_1
X_13916_ _06624_ _06204_ _06644_ _06639_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__o211a_1
X_17684_ _10160_ _10164_ _10193_ VGND VGND VPWR VPWR _10194_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_57_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14896_ _07559_ _07568_ _07566_ VGND VGND VPWR VPWR _07579_ sky130_fd_sc_hd__a21o_1
XFILLER_0_187_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16635_ _09185_ _09202_ _09204_ _09184_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19423_ _01227_ _01258_ _04870_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__o21a_1
XFILLER_0_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13847_ _06198_ _06214_ _06212_ VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__and3_1
XFILLER_0_175_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16566_ _09108_ _09140_ VGND VGND VPWR VPWR _09142_ sky130_fd_sc_hd__and2_1
X_19354_ _01189_ _01190_ _11726_ _11727_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_71_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13778_ net1052 _05788_ _06521_ _06446_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18305_ _10726_ _10771_ VGND VGND VPWR VPWR _10772_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15517_ _08149_ VGND VGND VPWR VPWR _08150_ sky130_fd_sc_hd__buf_4
X_12729_ _05537_ _05538_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__xor2_1
X_19285_ net247 VGND VGND VPWR VPWR _11687_ sky130_fd_sc_hd__buf_6
XFILLER_0_139_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16497_ _09072_ _09074_ VGND VGND VPWR VPWR _09075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18236_ _10656_ _10678_ _10704_ VGND VGND VPWR VPWR _10705_ sky130_fd_sc_hd__o21a_1
XFILLER_0_217_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15448_ _08051_ _08052_ _08089_ VGND VGND VPWR VPWR _08090_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_128_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18167_ _06701_ VGND VGND VPWR VPWR _10639_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15379_ _07949_ _07984_ VGND VGND VPWR VPWR _08023_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17118_ _09623_ _09668_ VGND VGND VPWR VPWR _09669_ sky130_fd_sc_hd__xor2_1
Xhold404 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[17\] VGND
+ VGND VPWR VPWR net586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18098_ top_inst.grid_inst.data_path_wires\[12\]\[3\] VGND VGND VPWR VPWR _10585_
+ sky130_fd_sc_hd__clkbuf_4
Xhold415 _00212_ VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 top_inst.deskew_buff_inst.col_input\[119\] VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold437 top_inst.axis_out_inst.out_buff_data\[96\] VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold448 top_inst.deskew_buff_inst.col_input\[122\] VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17049_ _09595_ _09600_ _09601_ VGND VGND VPWR VPWR _09602_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold459 _00023_ VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap178 net179 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20060_ _01873_ _01874_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23750_ clknet_leaf_135_clk net293 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20962_ _02695_ _02698_ _02729_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__nand3_1
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_205_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22701_ _04369_ _04373_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__xor2_2
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23681_ clknet_leaf_117_clk net438 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20893_ _02636_ _02662_ _02663_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__o21a_1
XFILLER_0_71_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22632_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[21\] _03937_ VGND
+ VGND VPWR VPWR _04308_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_193_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_1386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22563_ _04092_ _04241_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_499 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24302_ clknet_leaf_138_clk _00835_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[77\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21514_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[12\] _03080_ VGND
+ VGND VPWR VPWR _03247_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22494_ _04126_ _04147_ _04175_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24233_ clknet_leaf_112_clk _00766_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_181_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21445_ _03171_ _03179_ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_161_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24164_ clknet_leaf_9_clk _00697_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21376_ _03072_ _03112_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__xor2_1
XFILLER_0_160_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23115_ _04657_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__buf_4
XFILLER_0_47_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20327_ _02112_ _02113_ _02114_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__nand3_1
XFILLER_0_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24095_ clknet_leaf_99_clk _00628_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23046_ net3 _04615_ _04618_ _04619_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__o211a_1
X_20258_ net779 _01202_ _02047_ _02048_ _01863_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__o221a_1
XFILLER_0_101_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20189_ top_inst.grid_inst.data_path_wires\[16\]\[3\] VGND VGND VPWR VPWR _01995_
+ sky130_fd_sc_hd__buf_4
XFILLER_0_215_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_231_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14750_ _07398_ _07403_ net1124 VGND VGND VPWR VPWR _07438_ sky130_fd_sc_hd__a21oi_1
XTAP_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23948_ clknet_leaf_81_clk _00481_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11962_ net914 _04990_ _04992_ _04981_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__o211a_1
XTAP_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13701_ net1061 _05788_ _06445_ _06446_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__o211a_1
XTAP_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _07368_ _07369_ VGND VGND VPWR VPWR _07370_ sky130_fd_sc_hd__nor2_1
XFILLER_0_212_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23879_ clknet_leaf_61_clk _00412_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ net636 _04951_ _04953_ _04942_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16420_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[11\] VGND VGND
+ VPWR VPWR _08999_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13632_ _06377_ _06378_ VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__or2_1
X_16351_ top_inst.grid_inst.data_path_wires\[8\]\[7\] _08688_ VGND VGND VPWR VPWR
+ _08932_ sky130_fd_sc_hd__nand2_4
XFILLER_0_27_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13563_ _06273_ _06311_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_81_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15302_ _07947_ VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_212_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12514_ _05280_ _05279_ _05318_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__and3_1
XFILLER_0_183_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19070_ _11441_ _11448_ _11489_ VGND VGND VPWR VPWR _11490_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_152_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16282_ _08825_ _08827_ _08824_ VGND VGND VPWR VPWR _08865_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_164_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13494_ top_inst.grid_inst.data_path_wires\[2\]\[4\] top_inst.grid_inst.data_path_wires\[2\]\[3\]
+ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__nand4_1
XFILLER_0_136_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18021_ _10377_ _10502_ VGND VGND VPWR VPWR _10523_ sky130_fd_sc_hd__nor2_1
XFILLER_0_212_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15233_ _07877_ _07879_ VGND VGND VPWR VPWR _07880_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_858 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1018 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12445_ _05271_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_180_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15164_ _07774_ _07776_ _07773_ VGND VGND VPWR VPWR _07813_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_22_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12376_ net402 _05222_ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14115_ _06824_ _06787_ VGND VGND VPWR VPWR _06830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19972_ _01772_ _01773_ _01788_ _01789_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__o22a_1
X_15095_ top_inst.grid_inst.data_path_wires\[6\]\[0\] _07640_ _07637_ _07608_ VGND
+ VGND VPWR VPWR _07745_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_205_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14046_ _06758_ _06759_ _06761_ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__o21a_1
X_18923_ _11145_ _11154_ _11344_ _11345_ VGND VGND VPWR VPWR _11346_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_235_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18854_ _11277_ _11278_ VGND VGND VPWR VPWR _11279_ sky130_fd_sc_hd__nor2_1
XTAP_6470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17805_ _10310_ _10312_ VGND VGND VPWR VPWR _10313_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18785_ _11210_ _11211_ VGND VGND VPWR VPWR _11212_ sky130_fd_sc_hd__nand2_2
X_15997_ _08532_ _08604_ VGND VGND VPWR VPWR _08606_ sky130_fd_sc_hd__and2_1
XFILLER_0_237_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_238_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14948_ _04865_ _07378_ VGND VGND VPWR VPWR _07616_ sky130_fd_sc_hd__nand2_1
X_17736_ _10029_ _10054_ VGND VGND VPWR VPWR _10245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_221_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_221_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14879_ _07450_ _07562_ VGND VGND VPWR VPWR _07563_ sky130_fd_sc_hd__xor2_2
XFILLER_0_212_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17667_ _10166_ _10177_ VGND VGND VPWR VPWR _10178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_230_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19406_ _11701_ _11677_ _01240_ _01241_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__and4_1
X_16618_ _09185_ _09187_ _09190_ _09184_ VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17598_ _10089_ _10110_ VGND VGND VPWR VPWR _10111_ sky130_fd_sc_hd__xor2_2
XFILLER_0_106_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16549_ _09123_ _09124_ VGND VGND VPWR VPWR _09125_ sky130_fd_sc_hd__or2b_1
XFILLER_0_163_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19337_ _11729_ _11730_ VGND VGND VPWR VPWR _11731_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19268_ net985 _11662_ _11675_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18219_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[3\] _10686_ _10687_
+ VGND VGND VPWR VPWR _10688_ sky130_fd_sc_hd__a21bo_1
X_19199_ _11585_ _11615_ VGND VGND VPWR VPWR _11616_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21230_ _02966_ _02969_ VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__xor2_2
XFILLER_0_143_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold201 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[31\] VGND
+ VGND VPWR VPWR net383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[6\] VGND VGND
+ VPWR VPWR net394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 _00957_ VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold234 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[4\] VGND VGND
+ VPWR VPWR net416 sky130_fd_sc_hd__dlygate4sd3_1
X_21161_ _02902_ _02903_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[1\]
+ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__a21o_1
Xhold245 _00209_ VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold256 _00214_ VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[12\] VGND
+ VGND VPWR VPWR net449 sky130_fd_sc_hd__dlygate4sd3_1
X_20112_ _01899_ _01923_ _01914_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__nand3_1
Xhold278 top_inst.axis_out_inst.out_buff_data\[111\] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold289 top_inst.deskew_buff_inst.col_input\[126\] VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21092_ _02815_ _02842_ _02845_ _02846_ _02853_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__o221a_1
XFILLER_0_141_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_238_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20043_ _01857_ _01858_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23802_ clknet_leaf_77_clk _00335_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21994_ _03698_ _05275_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__or2_1
XFILLER_0_240_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 _05275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_217_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23733_ clknet_leaf_126_clk net457 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20945_ _02663_ _02708_ _02713_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_240_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23664_ clknet_leaf_132_clk net340 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20876_ _02473_ _02647_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22615_ _04290_ _04291_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__and2b_1
XFILLER_0_119_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23595_ clknet_leaf_100_clk _00128_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22546_ _04214_ _04224_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22477_ _04159_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24216_ clknet_leaf_19_clk _00749_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_12230_ net911 _05137_ _05146_ _05141_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__o211a_1
XFILLER_0_224_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21428_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[9\] _03122_ _03123_
+ VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24147_ clknet_leaf_16_clk _00680_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[13\]\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_20_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12161_ net373 _05097_ _05106_ _05101_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__o211a_1
X_21359_ _03093_ _03095_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__xor2_2
XFILLER_0_202_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12092_ net563 _05058_ _05067_ _05062_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__o211a_1
X_24078_ clknet_leaf_113_clk _00611_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold790 top_inst.axis_out_inst.out_buff_data\[31\] VGND VGND VPWR VPWR net972 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23029_ net27 _04601_ _04609_ _04606_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__o211a_1
XTAP_5010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15920_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[11\] _08452_ _08373_
+ VGND VGND VPWR VPWR _08531_ sky130_fd_sc_hd__a21o_1
XTAP_5021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15851_ _08421_ _08423_ VGND VGND VPWR VPWR _08464_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14802_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[13\] _07364_ VGND
+ VGND VPWR VPWR _07488_ sky130_fd_sc_hd__xnor2_1
XTAP_5098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18570_ _11005_ _11030_ VGND VGND VPWR VPWR _11031_ sky130_fd_sc_hd__xor2_1
X_15782_ _08349_ _08393_ VGND VGND VPWR VPWR _08396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_203_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ _05317_ _05779_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__nand2_1
XTAP_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14733_ _07419_ _07420_ VGND VGND VPWR VPWR _07421_ sky130_fd_sc_hd__nand2_1
X_17521_ _10044_ _09199_ VGND VGND VPWR VPWR _10045_ sky130_fd_sc_hd__or2_1
XTAP_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1056 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11945_ net1021 _04977_ _04983_ _04981_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _09931_ _09986_ _09968_ _09988_ _09967_ VGND VGND VPWR VPWR _09989_ sky130_fd_sc_hd__a32o_1
XFILLER_0_129_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _07350_ _07353_ VGND VGND VPWR VPWR _07354_ sky130_fd_sc_hd__xor2_4
XFILLER_0_86_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ net611 _04938_ _04944_ _04942_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__o211a_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16403_ _08937_ _08943_ _08982_ VGND VGND VPWR VPWR _08983_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13615_ _05886_ _06362_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__and2_1
X_17383_ _09901_ _09893_ VGND VGND VPWR VPWR _09923_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14595_ _07079_ _07078_ _07082_ _07074_ VGND VGND VPWR VPWR _07286_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_32_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16334_ _08914_ _08915_ VGND VGND VPWR VPWR _08916_ sky130_fd_sc_hd__and2_1
X_19122_ _11506_ _11507_ _11539_ VGND VGND VPWR VPWR _11541_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13546_ _06181_ _06214_ _06212_ _06184_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19053_ _11471_ _11472_ VGND VGND VPWR VPWR _11473_ sky130_fd_sc_hd__and2b_1
X_16265_ top_inst.grid_inst.data_path_wires\[8\]\[7\] _08676_ _08686_ _08682_ VGND
+ VGND VPWR VPWR _08848_ sky130_fd_sc_hd__nand4_1
XFILLER_0_36_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13477_ _06181_ _06208_ _06205_ _06184_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_113_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15216_ _07862_ _07863_ VGND VGND VPWR VPWR _07864_ sky130_fd_sc_hd__and2_1
X_18004_ _10497_ _10506_ VGND VGND VPWR VPWR _10507_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12428_ net680 _05256_ _05258_ _05247_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__o211a_1
XFILLER_0_242_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16196_ _08726_ _08746_ VGND VGND VPWR VPWR _08781_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15147_ top_inst.grid_inst.data_path_wires\[6\]\[7\] _07621_ _07629_ _07626_ VGND
+ VGND VPWR VPWR _07796_ sky130_fd_sc_hd__nand4_1
XFILLER_0_23_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12359_ net664 _05217_ _05219_ _05208_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19955_ _01759_ _01774_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__xnor2_1
X_15078_ _07710_ _07728_ VGND VGND VPWR VPWR _07729_ sky130_fd_sc_hd__xor2_2
XFILLER_0_227_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14029_ _06628_ _06643_ _06743_ _06744_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__nand4_1
X_18906_ _11328_ _11329_ VGND VGND VPWR VPWR _11330_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19886_ _01691_ _01708_ VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__xor2_1
XFILLER_0_177_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18837_ _11237_ _11245_ VGND VGND VPWR VPWR _11262_ sky130_fd_sc_hd__and2_1
XFILLER_0_222_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18768_ _11138_ _11135_ _11152_ _11149_ VGND VGND VPWR VPWR _11196_ sky130_fd_sc_hd__nand4_2
XFILLER_0_222_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17719_ _09661_ _10228_ VGND VGND VPWR VPWR _10229_ sky130_fd_sc_hd__and2_1
XFILLER_0_222_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18699_ _10606_ _10584_ _11141_ _11137_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_212_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20730_ _02506_ _02507_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20661_ _02366_ _02440_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22400_ _04083_ _04084_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__and2_1
X_23380_ net53 _04805_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__or2_1
X_20592_ _02363_ _02373_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22331_ _03695_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[2\] _03984_
+ _03983_ _03693_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__a32o_1
XFILLER_0_115_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_1290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22262_ top_inst.grid_inst.data_path_wires\[18\]\[7\] top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[2\]
+ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__nand2_4
XFILLER_0_115_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_1165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24001_ clknet_leaf_81_clk _00534_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21213_ _02951_ _02953_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__xor2_2
XFILLER_0_108_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22193_ _03880_ _03881_ _05353_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__a21o_1
X_21144_ _02871_ _02881_ _02892_ _02880_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__o211a_1
XFILLER_0_228_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21075_ _02825_ _02827_ _02837_ _05313_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__o31ai_2
X_20026_ _01824_ _01837_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__nand2_1
XFILLER_0_232_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21977_ _03686_ _02869_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__or2_1
Xrebuffer60 _11676_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer71 _09529_ VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__buf_2
XFILLER_0_16_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23716_ clknet_leaf_121_clk _00249_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20928_ _02667_ _02697_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23647_ clknet_leaf_127_clk _00180_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20859_ _02614_ _02631_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_166_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13400_ _06054_ _06150_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14380_ net1122 VGND VGND VPWR VPWR _07082_ sky130_fd_sc_hd__buf_2
XFILLER_0_147_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23578_ clknet_leaf_107_clk _00111_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13331_ _06104_ _06105_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22529_ _04208_ _04209_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16050_ _08651_ _08656_ VGND VGND VPWR VPWR _08657_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_228_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13262_ _06005_ _06002_ _06037_ _05405_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_150_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15001_ _07606_ _07631_ VGND VGND VPWR VPWR _07655_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12213_ net589 _05129_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__or2_1
X_13193_ _05744_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[6\] _05969_
+ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12144_ net835 _05084_ _05096_ _05088_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19740_ _01528_ _01567_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__xor2_2
X_16952_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[4\] net203 _09218_
+ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _09507_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12075_ net780 _05045_ _05057_ _05049_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__o211a_1
XFILLER_0_217_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15903_ _08476_ _08514_ _05335_ VGND VGND VPWR VPWR _08515_ sky130_fd_sc_hd__mux2_1
X_19671_ _01497_ _01498_ _01499_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16883_ _09436_ _09437_ _09438_ VGND VGND VPWR VPWR _09440_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18622_ _11079_ _11080_ VGND VGND VPWR VPWR _11081_ sky130_fd_sc_hd__nor2_1
XTAP_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15834_ _08409_ _08446_ VGND VGND VPWR VPWR _08447_ sky130_fd_sc_hd__xor2_1
XFILLER_0_235_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ _10591_ _10857_ _11013_ VGND VGND VPWR VPWR _11014_ sky130_fd_sc_hd__or3_1
XFILLER_0_235_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12977_ _05746_ _05756_ _05766_ _05767_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__o211a_1
XTAP_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15765_ _08370_ _08327_ _08378_ VGND VGND VPWR VPWR _08380_ sky130_fd_sc_hd__nor3_1
XFILLER_0_204_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17504_ _04865_ VGND VGND VPWR VPWR _10033_ sky130_fd_sc_hd__clkbuf_4
XTAP_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14716_ _07365_ _07370_ _07368_ VGND VGND VPWR VPWR _07404_ sky130_fd_sc_hd__a21o_1
X_11928_ net892 _04964_ _04973_ _04968_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15696_ top_inst.grid_inst.data_path_wires\[7\]\[0\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _08312_ sky130_fd_sc_hd__or2b_1
X_18484_ _10889_ _10905_ _10904_ VGND VGND VPWR VPWR _10947_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_234_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14647_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[5\] _07078_ _07334_
+ _07335_ VGND VGND VPWR VPWR _07337_ sky130_fd_sc_hd__a22o_1
X_17435_ _09935_ _09956_ _09954_ VGND VGND VPWR VPWR _09972_ sky130_fd_sc_hd__o21a_1
XFILLER_0_170_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11859_ net938 _04925_ _04934_ _04929_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_18 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_29 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14578_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[7\] _07269_ _06701_
+ VGND VGND VPWR VPWR _07270_ sky130_fd_sc_hd__mux2_1
X_17366_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[24\] _09494_ VGND
+ VGND VPWR VPWR _09907_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19105_ _11520_ _11522_ _11523_ VGND VGND VPWR VPWR _11524_ sky130_fd_sc_hd__nor3_1
XFILLER_0_15_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16317_ _08840_ _08842_ _08898_ VGND VGND VPWR VPWR _08899_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13529_ _06263_ _06278_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__xnor2_1
X_17297_ _09839_ _09840_ VGND VGND VPWR VPWR _09841_ sky130_fd_sc_hd__xor2_1
XFILLER_0_153_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19036_ _11428_ _11429_ _11456_ VGND VGND VPWR VPWR _11457_ sky130_fd_sc_hd__a21o_1
X_16248_ _04873_ VGND VGND VPWR VPWR _08831_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput103 net103 VGND VGND VPWR VPWR output_tdata[43] sky130_fd_sc_hd__clkbuf_4
X_16179_ _08695_ _08661_ VGND VGND VPWR VPWR _08764_ sky130_fd_sc_hd__nand2_1
Xoutput114 net114 VGND VGND VPWR VPWR output_tdata[53] sky130_fd_sc_hd__buf_2
Xoutput125 net125 VGND VGND VPWR VPWR output_tdata[63] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput136 net136 VGND VGND VPWR VPWR output_tdata[73] sky130_fd_sc_hd__clkbuf_4
Xoutput147 net147 VGND VGND VPWR VPWR output_tdata[83] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput158 net158 VGND VGND VPWR VPWR output_tdata[93] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_177_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19938_ _01736_ _01748_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__nand2_1
XFILLER_0_227_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19869_ _01691_ _01692_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__nor2_1
XFILLER_0_207_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21900_ _03453_ _03617_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__xnor2_1
X_22880_ _02706_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__buf_2
XFILLER_0_37_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21831_ _03516_ _03551_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__and2_1
XFILLER_0_218_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24550_ clknet_leaf_100_clk _01083_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dfxtp_2
X_21762_ _03469_ _03486_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23501_ clknet_leaf_140_clk _00034_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[91\]
+ sky130_fd_sc_hd__dfxtp_1
X_20713_ _06168_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__buf_4
X_24481_ clknet_leaf_46_clk _01014_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_valid
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_77_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21693_ _03405_ _03408_ _03407_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_93_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23432_ net817 _04827_ _04837_ _04831_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20644_ _02396_ _02401_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__and2_1
XFILLER_0_184_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23363_ net45 _04792_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20575_ _02004_ _02016_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[11\]
+ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22314_ _03945_ _03963_ _04000_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23294_ net139 _04753_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22245_ _03915_ _03917_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_239_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22176_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[5\] _03684_ VGND
+ VGND VPWR VPWR _03866_ sky130_fd_sc_hd__nand2_1
X_21127_ _02004_ _02877_ _02879_ _02880_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21058_ _02821_ _02822_ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__or2_1
XFILLER_0_233_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12900_ _05608_ _05704_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20009_ _01782_ _01825_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__nand2_1
X_13880_ _04862_ VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__buf_6
XFILLER_0_57_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_236_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12831_ _05601_ _05602_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__or2_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1064 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15550_ _08135_ _08155_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _08173_ sky130_fd_sc_hd__a21oi_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12762_ _05569_ _05570_ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__xnor2_2
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[6\] _07192_ _07193_
+ VGND VGND VPWR VPWR _07194_ sky130_fd_sc_hd__and3_1
XFILLER_0_185_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _08116_ _08118_ _08119_ _08121_ _05313_ VGND VGND VPWR VPWR _08122_ sky130_fd_sc_hd__o311a_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12693_ _05454_ _05459_ _05503_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__o21a_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17220_ _09748_ _09741_ _09763_ VGND VGND VPWR VPWR _09767_ sky130_fd_sc_hd__a21oi_1
X_14432_ _07126_ _07127_ VGND VGND VPWR VPWR _07128_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17151_ _09667_ _09669_ _09700_ VGND VGND VPWR VPWR _09701_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14363_ top_inst.skew_buff_inst.row\[1\].output_reg\[2\] top_inst.axis_in_inst.inbuf_bus\[10\]
+ net187 VGND VGND VPWR VPWR _07068_ sky130_fd_sc_hd__mux2_4
XFILLER_0_37_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput16 input_tdata[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_4
Xinput27 input_tdata[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_8
X_16102_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _08695_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13314_ _06086_ _06088_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_243_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17082_ _09630_ _09633_ VGND VGND VPWR VPWR _09634_ sky130_fd_sc_hd__xor2_2
X_14294_ _07002_ _07003_ VGND VGND VPWR VPWR _07004_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16033_ _08638_ _08639_ VGND VGND VPWR VPWR _08641_ sky130_fd_sc_hd__nand2_1
XFILLER_0_243_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13245_ _06020_ _06007_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__and2b_1
XFILLER_0_161_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13176_ _05901_ _05910_ _05954_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__o21a_1
XFILLER_0_236_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12127_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[27\] _05076_
+ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_1206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17984_ _10452_ _10456_ _10454_ VGND VGND VPWR VPWR _10487_ sky130_fd_sc_hd__a21o_1
XFILLER_0_236_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19723_ _01550_ _01551_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__or2_1
X_16935_ _09489_ _09490_ VGND VGND VPWR VPWR _09491_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_165_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12058_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[29\] _05036_
+ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__or2_1
XFILLER_0_236_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19654_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[3\]
+ _11708_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__and3_1
X_16866_ _09198_ _09215_ VGND VGND VPWR VPWR _09423_ sky130_fd_sc_hd__nand2_1
X_18605_ _11042_ _11064_ VGND VGND VPWR VPWR _11065_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_204_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15817_ _08429_ _08430_ VGND VGND VPWR VPWR _08431_ sky130_fd_sc_hd__or2_1
XFILLER_0_220_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19585_ _01362_ _01370_ _01369_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_137_1262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16797_ _09262_ _09289_ _09320_ _09355_ _09318_ VGND VGND VPWR VPWR _09356_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18536_ _10952_ _10997_ VGND VGND VPWR VPWR _10998_ sky130_fd_sc_hd__xnor2_1
X_15748_ _08149_ _08159_ _08361_ _08362_ VGND VGND VPWR VPWR _08363_ sky130_fd_sc_hd__a22o_1
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18467_ _10924_ _10929_ VGND VGND VPWR VPWR _10930_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15679_ _08293_ _08294_ _08295_ VGND VGND VPWR VPWR _08296_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17418_ _09954_ _09955_ VGND VGND VPWR VPWR _09956_ sky130_fd_sc_hd__nand2_2
XFILLER_0_157_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18398_ _10854_ _10862_ VGND VGND VPWR VPWR _10863_ sky130_fd_sc_hd__xor2_1
XFILLER_0_172_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17349_ _09826_ _09850_ _09851_ VGND VGND VPWR VPWR _09890_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1032 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20360_ _02145_ _02146_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19019_ _11145_ _11438_ _11439_ VGND VGND VPWR VPWR _11440_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20291_ _01989_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[3\] _02051_
+ _01992_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22030_ _03703_ _03680_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__nand2_1
XFILLER_0_228_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23981_ clknet_leaf_88_clk _00514_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_215_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22932_ net918 _04548_ _04553_ _04551_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22863_ net294 _04504_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24602_ clknet_leaf_23_clk _01135_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_39_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1069 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21814_ _03534_ _03535_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_210_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22794_ _04462_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24533_ clknet_leaf_130_clk _01066_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_78_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21745_ _03375_ _03452_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__nor2_1
XFILLER_0_210_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24464_ clknet_leaf_54_clk _00997_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21676_ _03375_ _03382_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__or2b_1
XFILLER_0_188_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23415_ top_inst.axis_out_inst.out_buff_data\[97\] _04596_ VGND VGND VPWR VPWR _04828_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_190_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20627_ _02366_ _02407_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__xnor2_1
X_24395_ clknet_leaf_37_clk _00928_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23346_ net164 _04779_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20558_ _02314_ _02340_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__xor2_2
XFILLER_0_225_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23277_ net131 _04740_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__or2_1
XFILLER_0_225_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20489_ _02236_ _02251_ _02252_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__and3_1
X_13030_ _05765_ _05811_ _05812_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__a21bo_1
X_22228_ _03859_ _03873_ _03916_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__o21a_1
XFILLER_0_218_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22159_ _03821_ _03830_ _03832_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_218_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_203_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14981_ _05755_ VGND VGND VPWR VPWR _07639_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_234_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16720_ _09278_ _09279_ _09273_ VGND VGND VPWR VPWR _09281_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13932_ _06637_ _06618_ _05328_ VGND VGND VPWR VPWR _06655_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_1272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16651_ top_inst.skew_buff_inst.row\[2\].output_reg\[7\] top_inst.axis_in_inst.inbuf_bus\[23\]
+ net185 VGND VGND VPWR VPWR _09217_ sky130_fd_sc_hd__mux2_2
X_13863_ _06602_ _06603_ VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12814_ _05579_ _05585_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15602_ _08219_ _08220_ VGND VGND VPWR VPWR _08221_ sky130_fd_sc_hd__nand2_1
X_19370_ _01185_ _01205_ _01206_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__or3_4
XFILLER_0_186_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16582_ _09151_ _09155_ VGND VGND VPWR VPWR _09157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13794_ _06535_ _06536_ VGND VGND VPWR VPWR _06537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18321_ _10754_ _10758_ VGND VGND VPWR VPWR _10787_ sky130_fd_sc_hd__nor2_1
X_12745_ _05552_ _05553_ _05509_ _05512_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__o211ai_4
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15533_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _08161_ sky130_fd_sc_hd__clkbuf_4
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15464_ _08005_ _08104_ VGND VGND VPWR VPWR _08105_ sky130_fd_sc_hd__xnor2_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ _10718_ _10719_ VGND VGND VPWR VPWR _10720_ sky130_fd_sc_hd__nand2_1
X_12676_ _05461_ _05470_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17203_ _09731_ _09733_ VGND VGND VPWR VPWR _09751_ sky130_fd_sc_hd__nand2_1
X_14415_ _07110_ _07111_ VGND VGND VPWR VPWR _07112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15395_ _07956_ _08037_ VGND VGND VPWR VPWR _08038_ sky130_fd_sc_hd__nand2_1
X_18183_ _10652_ _10653_ VGND VGND VPWR VPWR _10654_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_167_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17134_ _09630_ _09633_ _09684_ VGND VGND VPWR VPWR _09685_ sky130_fd_sc_hd__a21o_1
X_14346_ _07052_ _07053_ VGND VGND VPWR VPWR _07054_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold608 top_inst.deskew_buff_inst.col_input\[29\] VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__dlygate4sd3_1
X_17065_ _09616_ _09617_ VGND VGND VPWR VPWR _09618_ sky130_fd_sc_hd__nand2_1
XFILLER_0_204_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14277_ _06985_ _06986_ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__nand2_1
Xhold619 top_inst.axis_out_inst.out_buff_data\[124\] VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16016_ _08197_ _08624_ VGND VGND VPWR VPWR _08625_ sky130_fd_sc_hd__and2_1
X_13228_ _05998_ _06000_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13159_ _05750_ _05761_ _05935_ _05936_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__and4_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _10458_ _10428_ _10469_ VGND VGND VPWR VPWR _10471_ sky130_fd_sc_hd__nand3_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19706_ _01297_ _01314_ _11699_ _11704_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__or4b_4
X_16918_ _09471_ _09472_ _09470_ VGND VGND VPWR VPWR _09474_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17898_ _10354_ _10357_ VGND VGND VPWR VPWR _10403_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19637_ _01382_ _01383_ _01390_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_75_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16849_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[7\] _08066_ _09405_
+ _09406_ VGND VGND VPWR VPWR _09407_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19568_ _01398_ _01399_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18519_ _10979_ _10980_ VGND VGND VPWR VPWR _10981_ sky130_fd_sc_hd__nor2_1
XFILLER_0_220_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_929 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19499_ net241 _01331_ _01332_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__nor3_2
XFILLER_0_8_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21530_ _03210_ _03218_ _03262_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21461_ _02135_ _03195_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23200_ net94 _04701_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20412_ _02194_ _02195_ _02196_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__a21o_1
X_24180_ clknet_leaf_29_clk _00713_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21392_ _03126_ _03127_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23131_ net541 _04656_ _04667_ _04662_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20343_ _02127_ _02130_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23062_ net11 _04615_ _04627_ _04619_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__o211a_1
X_20274_ _02061_ _02062_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[3\]
+ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__o21bai_1
XTAP_6107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22013_ _03711_ _05275_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__or2_1
XTAP_6129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23964_ clknet_leaf_88_clk _00497_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22915_ _06619_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_242_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23895_ clknet_leaf_51_clk _00428_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22846_ _06619_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__buf_2
XFILLER_0_116_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_929 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22777_ _04390_ _04445_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__or2_1
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _05340_ _05344_ VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__or2_1
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24516_ clknet_leaf_133_clk _01049_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dfxtp_1
X_21728_ _03453_ _03428_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__nor2_1
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24447_ clknet_leaf_63_clk _00980_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[0\].output_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12461_ _05270_ _05283_ _05285_ _05261_ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21659_ _03348_ _03360_ _03359_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__a21oi_1
X_14200_ _06910_ _06912_ VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__xor2_1
X_15180_ _07826_ _07827_ VGND VGND VPWR VPWR _07828_ sky130_fd_sc_hd__xnor2_2
X_24378_ clknet_leaf_38_clk _00911_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12392_ net449 _05230_ _05238_ _05234_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14131_ _06842_ _06844_ _05633_ VGND VGND VPWR VPWR _06846_ sky130_fd_sc_hd__a21o_1
X_23329_ net156 _04779_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_205_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14062_ _06630_ _06643_ _06776_ _06777_ VGND VGND VPWR VPWR _06778_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13013_ _05791_ _05796_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18870_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[6\] _11294_ _08307_
+ VGND VGND VPWR VPWR _11295_ sky130_fd_sc_hd__mux2_1
XTAP_6630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17821_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[9\] _10236_ _10283_
+ VGND VGND VPWR VPWR _10328_ sky130_fd_sc_hd__a21o_1
XTAP_6663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17752_ _10258_ _10260_ VGND VGND VPWR VPWR _10261_ sky130_fd_sc_hd__xor2_1
XTAP_5973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14964_ _07627_ _07075_ VGND VGND VPWR VPWR _07628_ sky130_fd_sc_hd__or2_1
XTAP_5984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16703_ _08831_ _09264_ VGND VGND VPWR VPWR _09265_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13915_ _06643_ _06641_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17683_ _10159_ _10165_ VGND VGND VPWR VPWR _10193_ sky130_fd_sc_hd__or2b_1
XFILLER_0_215_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14895_ _07550_ _07552_ _07573_ VGND VGND VPWR VPWR _07578_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19422_ _01256_ _01257_ _06168_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__and3b_1
X_16634_ _09203_ _09199_ VGND VGND VPWR VPWR _09204_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13846_ _06541_ _06570_ _06586_ VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__o21a_1
XFILLER_0_186_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19353_ _11726_ _11727_ _01189_ _01190_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_130_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16565_ _09108_ _09140_ VGND VGND VPWR VPWR _09141_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13777_ _06519_ _06520_ _05328_ VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18304_ _10767_ _10770_ VGND VGND VPWR VPWR _10771_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15516_ top_inst.grid_inst.data_path_wires\[7\]\[6\] VGND VGND VPWR VPWR _08149_
+ sky130_fd_sc_hd__buf_2
X_19284_ top_inst.skew_buff_inst.row\[3\].output_reg\[2\] top_inst.axis_in_inst.inbuf_bus\[26\]
+ net188 VGND VGND VPWR VPWR _11686_ sky130_fd_sc_hd__mux2_4
X_12728_ _05284_ _05306_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__nand2_2
XFILLER_0_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_927 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16496_ _09035_ _09036_ _09073_ VGND VGND VPWR VPWR _09074_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18235_ _10675_ _10677_ VGND VGND VPWR VPWR _10704_ sky130_fd_sc_hd__or2b_1
X_12659_ _05461_ _05470_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15447_ _08053_ _08054_ VGND VGND VPWR VPWR _08089_ sky130_fd_sc_hd__or2b_1
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18166_ _10626_ _10637_ VGND VGND VPWR VPWR _10638_ sky130_fd_sc_hd__xnor2_1
X_15378_ _07982_ _08021_ VGND VGND VPWR VPWR _08022_ sky130_fd_sc_hd__xor2_2
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17117_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[14\] _09419_ VGND
+ VGND VPWR VPWR _09668_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14329_ _07036_ _07037_ VGND VGND VPWR VPWR _07038_ sky130_fd_sc_hd__nor2_1
Xhold405 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[15\] VGND
+ VGND VPWR VPWR net587 sky130_fd_sc_hd__dlygate4sd3_1
X_18097_ _10583_ VGND VGND VPWR VPWR _10584_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold416 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[29\] VGND
+ VGND VPWR VPWR net598 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold427 _01176_ VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold438 top_inst.valid_pipe\[7\] VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__dlygate4sd3_1
X_17048_ _09598_ _09599_ _09597_ VGND VGND VPWR VPWR _09601_ sky130_fd_sc_hd__a21o_1
Xhold449 top_inst.deskew_buff_inst.col_input\[42\] VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap168 _01790_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap179 _02233_ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18999_ _11417_ _11419_ VGND VGND VPWR VPWR _11421_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20961_ _02695_ _02698_ _02729_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__a21o_1
XFILLER_0_224_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22700_ _04371_ _04372_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__and2b_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23680_ clknet_leaf_117_clk net484 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20892_ _02629_ _02640_ _02658_ VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22631_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[20\] _04163_ _03938_
+ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22562_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[18\] _04163_ VGND
+ VGND VPWR VPWR _04241_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24301_ clknet_leaf_138_clk _00834_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[76\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21513_ _03245_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__clkbuf_4
X_22493_ _04146_ _04145_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__and2b_1
XFILLER_0_111_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_1141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24232_ clknet_leaf_111_clk _00765_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[16\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21444_ _03176_ _03178_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__xor2_2
XFILLER_0_32_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24163_ clknet_leaf_9_clk _00696_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_21375_ _03109_ _03111_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__xor2_2
XFILLER_0_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23114_ top_inst.axis_out_inst.out_buff_enabled _04857_ VGND VGND VPWR VPWR _04657_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_43_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20326_ _02078_ _02080_ _02079_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__a21bo_1
X_24094_ clknet_leaf_99_clk _00627_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23045_ _04550_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20257_ _02030_ _02036_ _02046_ _01984_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__a31o_1
XTAP_5203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20188_ _01993_ _10033_ _01994_ _01840_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__o211a_1
XTAP_5247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ top_inst.axis_out_inst.out_buff_data\[52\] _04982_ VGND VGND VPWR VPWR _04992_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_93_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23947_ clknet_leaf_85_clk _00480_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _05260_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__clkbuf_4
XTAP_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ _07367_ _07366_ VGND VGND VPWR VPWR _07369_ sky130_fd_sc_hd__and2b_1
XTAP_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23878_ clknet_leaf_51_clk _00411_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11892_ net474 _04943_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13631_ _06195_ _06205_ _06375_ _06376_ VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__and4_1
XFILLER_0_211_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22829_ _09787_ _04493_ _04494_ _03929_ VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16350_ _08928_ _08930_ VGND VGND VPWR VPWR _08931_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13562_ _06309_ _06310_ VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12513_ _05273_ _05283_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15301_ _07117_ _07946_ VGND VGND VPWR VPWR _07947_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16281_ _08822_ _08863_ VGND VGND VPWR VPWR _08864_ sky130_fd_sc_hd__xor2_1
XFILLER_0_136_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13493_ _06232_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18020_ _10413_ _10493_ _10495_ VGND VGND VPWR VPWR _10522_ sky130_fd_sc_hd__o21ai_1
X_12444_ top_inst.skew_buff_inst.row\[0\].output_reg\[0\] top_inst.axis_in_inst.inbuf_bus\[0\]
+ net211 VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__mux2_2
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15232_ _07878_ VGND VGND VPWR VPWR _07879_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15163_ _07771_ _07811_ VGND VGND VPWR VPWR _07812_ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12375_ net452 _05217_ _05228_ _05221_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14114_ _06824_ _06787_ _06827_ _06828_ VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19971_ _01772_ _01773_ _01788_ _01789_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__nor4_1
X_15094_ _07720_ _07726_ VGND VGND VPWR VPWR _07744_ sky130_fd_sc_hd__or2b_1
XFILLER_0_205_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14045_ _06758_ _06759_ _06761_ VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__nor3_1
X_18922_ _11143_ _11158_ _11140_ _11156_ VGND VGND VPWR VPWR _11345_ sky130_fd_sc_hd__nand4_2
XFILLER_0_201_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18853_ _11140_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[2\] _11275_
+ _11276_ VGND VGND VPWR VPWR _11278_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_235_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17804_ _10239_ _10257_ _10311_ VGND VGND VPWR VPWR _10312_ sky130_fd_sc_hd__a21oi_1
XTAP_6493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18784_ _11140_ _11138_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _11211_ sky130_fd_sc_hd__nand4_1
XTAP_5770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15996_ _08532_ _08604_ VGND VGND VPWR VPWR _08605_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17735_ _10242_ _10243_ VGND VGND VPWR VPWR _10244_ sky130_fd_sc_hd__nand2_1
XFILLER_0_206_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14947_ top_inst.grid_inst.data_path_wires\[6\]\[4\] VGND VGND VPWR VPWR _07615_
+ sky130_fd_sc_hd__buf_4
XFILLER_0_37_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_221_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17666_ _10167_ _10176_ VGND VGND VPWR VPWR _10177_ sky130_fd_sc_hd__xor2_1
X_14878_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[15\] _07364_ VGND
+ VGND VPWR VPWR _07562_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_216_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19405_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[2\] _11692_ _01238_
+ _01239_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16617_ _09189_ _08684_ VGND VGND VPWR VPWR _09190_ sky130_fd_sc_hd__or2_1
X_13829_ _06542_ _06570_ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_230_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17597_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[4\] _10109_ VGND
+ VGND VPWR VPWR _10110_ sky130_fd_sc_hd__xor2_2
XFILLER_0_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19336_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[1\] _11715_ _11716_
+ VGND VGND VPWR VPWR _11730_ sky130_fd_sc_hd__a21boi_1
X_16548_ _09117_ _09088_ _09122_ VGND VGND VPWR VPWR _09124_ sky130_fd_sc_hd__nand3_1
XFILLER_0_169_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_910 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19267_ net962 _11662_ _11675_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__o21a_1
X_16479_ _09055_ _09056_ VGND VGND VPWR VPWR _09057_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18218_ top_inst.grid_inst.data_path_wires\[12\]\[1\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[12\]\[2\]
+ VGND VGND VPWR VPWR _10687_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19198_ _11578_ _11614_ VGND VGND VPWR VPWR _11615_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_143_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18149_ _10599_ _10577_ _10600_ _10597_ VGND VGND VPWR VPWR _10622_ sky130_fd_sc_hd__nand4_2
XFILLER_0_108_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold202 _00198_ VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 _00908_ VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[3\] VGND VGND
+ VPWR VPWR net406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 _00938_ VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21160_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[1\] _02902_ _02903_
+ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__nand3_1
XFILLER_0_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold246 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[31\] VGND
+ VGND VPWR VPWR net428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold257 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[12\] VGND
+ VGND VPWR VPWR net439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20111_ _01899_ _01914_ _01923_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__a21o_1
Xhold268 _00275_ VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 top_inst.axis_out_inst.out_buff_data\[104\] VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21091_ _02819_ _02843_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__or2b_1
XFILLER_0_223_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20042_ _01855_ _01856_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__and2_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23801_ clknet_leaf_72_clk _00334_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21993_ _03697_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__clkbuf_4
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23732_ clknet_leaf_125_clk _00265_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_108 _05275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20944_ _02678_ _02685_ _02702_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__o21ai_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_119 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23663_ clknet_leaf_132_clk net376 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20875_ _02645_ _02646_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22614_ _04218_ _04289_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23594_ clknet_leaf_101_clk _00127_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22545_ _04214_ _04224_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_142_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_142_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22476_ _07707_ _04158_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24215_ clknet_leaf_118_clk _00748_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_21427_ _03125_ _03126_ _03127_ _03129_ _03124_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__a32o_1
XFILLER_0_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24146_ clknet_leaf_16_clk _00679_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[13\]\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_12160_ top_inst.axis_out_inst.out_buff_data\[9\] _05102_ VGND VGND VPWR VPWR _05106_
+ sky130_fd_sc_hd__or2_1
X_21358_ _02866_ _02893_ _03053_ _03094_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20309_ _02070_ _02096_ _02097_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__o21a_1
X_12091_ net1104 _05063_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__or2_1
X_24077_ clknet_leaf_113_clk _00610_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold780 top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[23\] VGND VGND
+ VPWR VPWR net962 sky130_fd_sc_hd__dlygate4sd3_1
X_21289_ _03026_ _03027_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold791 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[26\] VGND
+ VGND VPWR VPWR net973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23028_ top_inst.axis_in_inst.inbuf_bus\[4\] _04603_ VGND VGND VPWR VPWR _04609_
+ sky130_fd_sc_hd__or2_1
XTAP_5000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15850_ _08461_ _08462_ VGND VGND VPWR VPWR _08463_ sky130_fd_sc_hd__xnor2_1
XTAP_5066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_232_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[12\] _07364_ _07280_
+ VGND VGND VPWR VPWR _07487_ sky130_fd_sc_hd__a21o_1
XTAP_5088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _06848_ _08394_ _08395_ _08166_ VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__o211a_1
XTAP_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _05775_ _05777_ _05778_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__o21ai_1
XTAP_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _10044_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14732_ _07083_ _07086_ _07417_ _07418_ VGND VGND VPWR VPWR _07420_ sky130_fd_sc_hd__a22o_1
XTAP_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ net513 _04982_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__or2_1
XTAP_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17451_ _09951_ _09946_ VGND VGND VPWR VPWR _09988_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14663_ _07351_ _07352_ VGND VGND VPWR VPWR _07353_ sky130_fd_sc_hd__nand2_2
XFILLER_0_129_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11875_ net570 _04943_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__or2_1
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16402_ _08936_ _08934_ VGND VGND VPWR VPWR _08982_ sky130_fd_sc_hd__and2b_1
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13614_ _05887_ _06359_ _06360_ _06361_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__a31o_1
X_17382_ _09911_ _09921_ VGND VGND VPWR VPWR _09922_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14594_ _07070_ _07086_ VGND VGND VPWR VPWR _07285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19121_ _11506_ _11507_ _11539_ VGND VGND VPWR VPWR _11540_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16333_ _08873_ _08874_ _08913_ VGND VGND VPWR VPWR _08915_ sky130_fd_sc_hd__nand3_1
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13545_ _06264_ _06269_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__or2_1
XFILLER_0_171_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_133_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_133_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19052_ _11147_ _11154_ _11439_ _11438_ _11145_ VGND VGND VPWR VPWR _11472_ sky130_fd_sc_hd__a32o_1
XFILLER_0_180_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16264_ _08676_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[1\] _08682_
+ top_inst.grid_inst.data_path_wires\[8\]\[7\] VGND VGND VPWR VPWR _08847_ sky130_fd_sc_hd__a22o_1
X_13476_ net1056 _05788_ _06228_ _06207_ VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1011 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18003_ _10504_ _10505_ VGND VGND VPWR VPWR _10506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_1153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15215_ _07821_ _07822_ _07861_ VGND VGND VPWR VPWR _07863_ sky130_fd_sc_hd__nand3_1
X_12427_ net308 _05248_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__or2_1
X_16195_ _08763_ _08779_ VGND VGND VPWR VPWR _08780_ sky130_fd_sc_hd__xor2_1
XFILLER_0_112_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15146_ _07621_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[1\] _07626_
+ top_inst.grid_inst.data_path_wires\[6\]\[7\] VGND VGND VPWR VPWR _07795_ sky130_fd_sc_hd__a22o_1
X_12358_ net335 _05209_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19954_ _01772_ _01773_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__xor2_1
X_15077_ _07719_ _07727_ VGND VGND VPWR VPWR _07728_ sky130_fd_sc_hd__xor2_2
X_12289_ net495 _05169_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14028_ _06628_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[2\] _06743_
+ _06744_ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__a22o_1
X_18905_ _11291_ _11293_ _11290_ VGND VGND VPWR VPWR _11329_ sky130_fd_sc_hd__o21bai_2
X_19885_ _01704_ _01707_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_219_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18836_ _11238_ _11244_ VGND VGND VPWR VPWR _11261_ sky130_fd_sc_hd__or2b_1
XTAP_6290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18767_ _11135_ _11152_ _11149_ _11138_ VGND VGND VPWR VPWR _11195_ sky130_fd_sc_hd__a22o_1
X_15979_ _08509_ _08548_ VGND VGND VPWR VPWR _08589_ sky130_fd_sc_hd__and2b_1
XFILLER_0_222_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17718_ _10226_ _10227_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[7\]
+ _07816_ VGND VGND VPWR VPWR _10228_ sky130_fd_sc_hd__a2bb2o_1
X_18698_ _11140_ _11133_ VGND VGND VPWR VPWR _11141_ sky130_fd_sc_hd__or2_1
XFILLER_0_194_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17649_ _10050_ _10129_ _10131_ _10128_ VGND VGND VPWR VPWR _10160_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_37_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_808 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20660_ _02406_ _02439_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19319_ net917 _10616_ _11713_ _11714_ VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_124_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_124_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20591_ _02371_ _02372_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22330_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[10\] _03894_ _03938_
+ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22261_ _03946_ _03948_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24000_ clknet_leaf_83_clk _00533_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_182_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21212_ _02891_ _02925_ _02952_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__a21bo_1
X_22192_ _03880_ _03881_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21143_ _02891_ _02021_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21074_ _02825_ net228 _02837_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20025_ _01813_ _01836_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__nand2_1
XFILLER_0_225_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_1377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21976_ top_inst.grid_inst.data_path_wires\[18\]\[3\] VGND VGND VPWR VPWR _03686_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_240_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer50 _01266_ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer61 net242 VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_139_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer72 _09191_ VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__buf_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20927_ _02695_ _02696_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__nand2_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23715_ clknet_leaf_121_clk _00248_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20858_ _02629_ _02630_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__nand2_1
X_23646_ clknet_leaf_127_clk _00179_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_115_clk clknet_4_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23577_ clknet_leaf_107_clk _00110_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20789_ _02532_ _02564_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__xor2_1
XFILLER_0_107_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13330_ _06025_ _06072_ _06070_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__a21oi_1
X_22528_ _04177_ _04207_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13261_ _06005_ _06002_ _06037_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22459_ _04139_ _04140_ _04025_ _04136_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15000_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[1\] _06660_ _07654_
+ _07643_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__o211a_1
X_12212_ net383 _05123_ _05135_ _05128_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__o211a_1
X_13192_ _05744_ _05770_ _05969_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12143_ net677 _05089_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__or2_1
X_24129_ clknet_leaf_119_clk _00662_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16951_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[3\] net203 _09218_
+ VGND VGND VPWR VPWR _09506_ sky130_fd_sc_hd__and3_1
X_12074_ net558 _05050_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15902_ _08512_ _08513_ VGND VGND VPWR VPWR _08514_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_218_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19670_ _01497_ _01498_ _01499_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__nand3_2
XFILLER_0_159_1146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16882_ _09436_ _09437_ _09438_ VGND VGND VPWR VPWR _09439_ sky130_fd_sc_hd__nand3_2
XFILLER_0_216_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18621_ _10969_ _11078_ VGND VGND VPWR VPWR _11080_ sky130_fd_sc_hd__and2_1
XTAP_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15833_ _08150_ _08444_ _08445_ VGND VGND VPWR VPWR _08446_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_205_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18552_ top_inst.grid_inst.data_path_wires\[12\]\[7\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _11013_ sky130_fd_sc_hd__nand2_1
XFILLER_0_220_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _08370_ _08327_ _08378_ VGND VGND VPWR VPWR _08379_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12976_ _05260_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__clkbuf_4
XTAP_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17503_ top_inst.grid_inst.data_path_wires\[11\]\[4\] VGND VGND VPWR VPWR _10032_
+ sky130_fd_sc_hd__clkbuf_4
XTAP_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _07359_ _07400_ VGND VGND VPWR VPWR _07403_ sky130_fd_sc_hd__or2b_1
XTAP_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11927_ net676 _04969_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__or2_1
X_18483_ _10930_ _10945_ VGND VGND VPWR VPWR _10946_ sky130_fd_sc_hd__xor2_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15695_ top_inst.grid_inst.data_path_wires\[7\]\[1\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _08311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_213_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _09787_ _09969_ _09970_ _09971_ _09806_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__o311a_1
X_14646_ _07083_ _07078_ _07334_ _07335_ VGND VGND VPWR VPWR _07336_ sky130_fd_sc_hd__nand4_1
XFILLER_0_28_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ net337 _04930_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17365_ net252 _09905_ VGND VGND VPWR VPWR _09906_ sky130_fd_sc_hd__xor2_1
XFILLER_0_28_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_19 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_106_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_16
X_14577_ _07267_ _07268_ VGND VGND VPWR VPWR _07269_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11789_ net367 _04885_ _04894_ _04889_ VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19104_ _11164_ _11145_ _11521_ VGND VGND VPWR VPWR _11523_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16316_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[8\] _08897_ VGND
+ VGND VPWR VPWR _08898_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13528_ _06270_ _06277_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__xor2_2
X_17296_ _09726_ _09816_ VGND VGND VPWR VPWR _09840_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19035_ _11430_ _11455_ VGND VGND VPWR VPWR _11456_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16247_ _08830_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13459_ _06196_ _06204_ _06215_ _06207_ VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput104 net104 VGND VGND VPWR VPWR output_tdata[44] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16178_ _08749_ _08754_ VGND VGND VPWR VPWR _08763_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput115 net115 VGND VGND VPWR VPWR output_tdata[54] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput126 net126 VGND VGND VPWR VPWR output_tdata[64] sky130_fd_sc_hd__clkbuf_4
Xoutput137 net137 VGND VGND VPWR VPWR output_tdata[74] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15129_ _07117_ _07778_ VGND VGND VPWR VPWR _07779_ sky130_fd_sc_hd__and2_1
Xoutput148 net148 VGND VGND VPWR VPWR output_tdata[84] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput159 net159 VGND VGND VPWR VPWR output_tdata[94] sky130_fd_sc_hd__buf_2
XFILLER_0_227_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19937_ net925 _01735_ _01757_ _11714_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19868_ _01679_ _01680_ _01690_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_207_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18819_ _11238_ _11244_ VGND VGND VPWR VPWR _11245_ sky130_fd_sc_hd__xnor2_2
X_19799_ _01625_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21830_ _03375_ _03534_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__nor2_1
XFILLER_0_223_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21761_ _03484_ _03485_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__and2_1
XFILLER_0_194_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23500_ clknet_leaf_139_clk _00033_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[90\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20712_ _02490_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24480_ clknet_leaf_55_clk _01013_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21692_ net891 _06169_ _03419_ _02909_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23431_ net461 _04835_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__or2_1
XFILLER_0_190_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20643_ _02389_ _02419_ _02422_ VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_11_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23362_ net697 _04791_ _04799_ _04795_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20574_ _01997_ _02227_ _02325_ _02326_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_18_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22313_ _03960_ _03962_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23293_ net727 _04752_ _04760_ _04756_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__o211a_1
XFILLER_0_225_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22244_ _03919_ _03922_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__or2_2
XFILLER_0_225_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22175_ _03863_ _03864_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21126_ _02706_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21057_ _02794_ _02796_ _02820_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__and3_1
XFILLER_0_195_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20008_ _01783_ _01806_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_241_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12830_ _05613_ _05611_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__and2b_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _05298_ _05297_ VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__nand2_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21959_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[25\] _03672_ _03078_
+ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__a21o_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[0\]
+ _07081_ _07085_ VGND VGND VPWR VPWR _07193_ sky130_fd_sc_hd__nand4_1
XFILLER_0_189_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _05414_ _05453_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__or2_1
X_15480_ _08094_ _08095_ _08120_ _08092_ VGND VGND VPWR VPWR _08121_ sky130_fd_sc_hd__a211o_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14431_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[3\] _07070_ _07060_
+ _07065_ VGND VGND VPWR VPWR _07127_ sky130_fd_sc_hd__nand4_2
XFILLER_0_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23629_ clknet_leaf_102_clk net257 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17150_ _09625_ _09668_ VGND VGND VPWR VPWR _09700_ sky130_fd_sc_hd__nor2_1
X_14362_ _05290_ _07065_ _07067_ _06684_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput17 input_tdata[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_107_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16101_ _08671_ _08681_ _08694_ _08692_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__o211a_1
Xinput28 input_tdata[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_2
XFILLER_0_91_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13313_ _05753_ _05768_ _06087_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__and3_1
X_17081_ _09623_ _09632_ VGND VGND VPWR VPWR _09633_ sky130_fd_sc_hd__xor2_2
X_14293_ _06965_ _06969_ _07001_ VGND VGND VPWR VPWR _07003_ sky130_fd_sc_hd__or3_1
XFILLER_0_122_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13244_ _06007_ _06020_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__and2b_1
X_16032_ _08638_ _08639_ VGND VGND VPWR VPWR _08640_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_1000 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13175_ _05888_ _05900_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12126_ net274 _05084_ _05086_ _05075_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17983_ _10404_ _10442_ _10482_ _10485_ _10481_ VGND VGND VPWR VPWR _10486_ sky130_fd_sc_hd__a32o_1
XFILLER_0_97_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19722_ _01548_ _01549_ _01522_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__a21oi_1
X_16934_ _09413_ _09445_ _09443_ VGND VGND VPWR VPWR _09490_ sky130_fd_sc_hd__a21o_1
X_12057_ net869 _05045_ _05047_ _05035_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19653_ _01478_ _01482_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__xor2_1
X_16865_ _09414_ _09421_ VGND VGND VPWR VPWR _09422_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18604_ _11062_ _11063_ VGND VGND VPWR VPWR _11064_ sky130_fd_sc_hd__nand2_1
X_15816_ _08426_ _08428_ VGND VGND VPWR VPWR _08430_ sky130_fd_sc_hd__and2_1
X_19584_ _01413_ _01414_ _01406_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__a21o_1
XFILLER_0_204_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16796_ _09259_ _09289_ VGND VGND VPWR VPWR _09355_ sky130_fd_sc_hd__or2_1
XFILLER_0_220_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_467 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18535_ _10995_ _10996_ VGND VGND VPWR VPWR _10997_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_1176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15747_ _08147_ _08163_ _08164_ _08161_ VGND VGND VPWR VPWR _08362_ sky130_fd_sc_hd__nand4_4
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _05753_ _05735_ _05754_ _05743_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__o211a_1
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18466_ _10927_ _10928_ VGND VGND VPWR VPWR _10929_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15678_ _08247_ _08255_ VGND VGND VPWR VPWR _08295_ sky130_fd_sc_hd__and2_1
XFILLER_0_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17417_ _09625_ _09953_ VGND VGND VPWR VPWR _09955_ sky130_fd_sc_hd__nand2_1
X_14629_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[8\] _07281_ _07280_
+ VGND VGND VPWR VPWR _07319_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18397_ _10860_ _10861_ VGND VGND VPWR VPWR _10862_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17348_ _09867_ _09862_ VGND VGND VPWR VPWR _09889_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17279_ _09768_ _09823_ VGND VGND VPWR VPWR _09824_ sky130_fd_sc_hd__or2b_2
XFILLER_0_130_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19018_ top_inst.grid_inst.data_path_wires\[13\]\[6\] _11158_ _11156_ top_inst.grid_inst.data_path_wires\[13\]\[7\]
+ VGND VGND VPWR VPWR _11439_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20290_ _01992_ _01989_ _02013_ _02011_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__nand4_1
XFILLER_0_24_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_1109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_1319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23980_ clknet_leaf_87_clk _00513_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_243_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22931_ net704 _04543_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_719 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22862_ net986 _04509_ _04513_ _04511_ VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24601_ clknet_leaf_24_clk _01134_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_6_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21813_ _03375_ _03516_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__nor2_1
X_22793_ _04438_ _04456_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24532_ clknet_leaf_103_clk _01065_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_66_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21744_ _03399_ _03439_ _03466_ _03468_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_93_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24463_ clknet_leaf_59_clk _00996_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_21675_ _03377_ _03381_ _03379_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__a21o_1
XFILLER_0_171_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23414_ _05736_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__clkbuf_4
X_20626_ _02405_ _02406_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__xor2_1
X_24394_ clknet_leaf_38_clk _00927_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23345_ net575 _04778_ _04789_ _04782_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__o211a_1
X_20557_ _02338_ _02339_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23276_ net940 _04739_ _04750_ _04743_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20488_ _02251_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__inv_2
XFILLER_0_225_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22227_ _03860_ _03872_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__nand2_1
X_22158_ _03813_ _03818_ _03847_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_160_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21109_ _01993_ _11142_ _02867_ _02707_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__o211a_1
X_14980_ _07619_ _06647_ _07638_ _07618_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__o211a_1
X_22089_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[18\]\[2\]
+ top_inst.grid_inst.data_path_wires\[18\]\[1\] _03707_ VGND VGND VPWR VPWR _03781_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_238_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13931_ _06635_ _06647_ _06654_ _06639_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16650_ _09213_ _05276_ _09216_ _09184_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13862_ _06600_ _06601_ VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15601_ _08163_ top_inst.grid_inst.data_path_wires\[7\]\[3\] _08157_ _08154_ VGND
+ VGND VPWR VPWR _08220_ sky130_fd_sc_hd__nand4_1
X_12813_ _05619_ _05620_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__or2_1
XFILLER_0_241_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16581_ _09151_ _09155_ VGND VGND VPWR VPWR _09156_ sky130_fd_sc_hd__or2_1
X_13793_ _06523_ _06498_ _06534_ VGND VGND VPWR VPWR _06536_ sky130_fd_sc_hd__nand3_1
XFILLER_0_202_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18320_ _10786_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__clkbuf_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15532_ _08139_ _07639_ _08160_ _08142_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_1302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12744_ _05509_ _05512_ _05552_ _05553_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__a211o_2
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _10591_ top_inst.grid_inst.data_path_wires\[12\]\[5\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _10719_ sky130_fd_sc_hd__nand4_1
X_15463_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[15\] _07924_ VGND
+ VGND VPWR VPWR _08104_ sky130_fd_sc_hd__xnor2_2
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _05446_ _05460_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17202_ _09738_ _09725_ VGND VGND VPWR VPWR _09750_ sky130_fd_sc_hd__or2b_1
XFILLER_0_182_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14414_ _07070_ _07061_ _07109_ VGND VGND VPWR VPWR _07111_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18182_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[2\] _10629_ _10630_
+ VGND VGND VPWR VPWR _10653_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_37_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15394_ _08035_ _08036_ VGND VGND VPWR VPWR _08037_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17133_ _09625_ _09632_ VGND VGND VPWR VPWR _09684_ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_838 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14345_ _06981_ _07034_ _07032_ VGND VGND VPWR VPWR _07053_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17064_ _09584_ _09615_ VGND VGND VPWR VPWR _09617_ sky130_fd_sc_hd__nand2_1
Xhold609 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[25\] VGND
+ VGND VPWR VPWR net791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14276_ _06985_ _06986_ VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16015_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[14\] _08066_ _08622_
+ _08623_ VGND VGND VPWR VPWR _08624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13227_ net1024 _05788_ _06004_ _05767_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13158_ _05750_ _05761_ _05935_ _05936_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_236_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ net486 _05071_ _05077_ _05075_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13089_ _05868_ _05869_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__nor2_1
X_17966_ _10458_ _10428_ _10469_ VGND VGND VPWR VPWR _10470_ sky130_fd_sc_hd__a21o_1
XFILLER_0_236_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16917_ _09470_ _09471_ _09472_ VGND VGND VPWR VPWR _09473_ sky130_fd_sc_hd__nand3_1
X_19705_ _01533_ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17897_ net1038 _10364_ _10401_ _10402_ _09886_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__o221a_1
XFILLER_0_192_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16848_ _09403_ _09404_ _05399_ VGND VGND VPWR VPWR _09406_ sky130_fd_sc_hd__a21oi_1
X_19636_ _01432_ _01466_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_215_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19567_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[9\] _01354_ VGND
+ VGND VPWR VPWR _01399_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_215_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16779_ _09213_ _09211_ _09186_ _09192_ VGND VGND VPWR VPWR _09338_ sky130_fd_sc_hd__and4_1
X_18518_ _10977_ _10978_ _10975_ VGND VGND VPWR VPWR _10980_ sky130_fd_sc_hd__o21a_1
X_19498_ _01283_ _01285_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__and2b_1
XFILLER_0_48_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_662 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18449_ _10911_ _10912_ VGND VGND VPWR VPWR _10913_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21460_ top_inst.deskew_buff_inst.col_input\[74\] _05731_ _03193_ _03194_ VGND VGND
+ VPWR VPWR _03195_ sky130_fd_sc_hd__a22o_1
XFILLER_0_185_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20411_ _02194_ _02195_ _02196_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__nand3_1
XFILLER_0_16_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21391_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[9\] _03080_ VGND
+ VGND VPWR VPWR _03127_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_6__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_4_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23130_ net132 _04659_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20342_ _02066_ _02128_ _02129_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_222_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23061_ net1111 _04616_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20273_ _02061_ _02062_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[3\]
+ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__or3b_1
XFILLER_0_101_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22012_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _03711_ sky130_fd_sc_hd__buf_2
XTAP_6119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_228_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23963_ clknet_leaf_88_clk _00496_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_95_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_224_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22914_ net416 _04535_ _04542_ _04537_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23894_ clknet_leaf_51_clk _00427_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22845_ net394 _04496_ _04503_ _04498_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22776_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[27\] _04215_ _04216_
+ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__a21oi_2
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_969 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24515_ clknet_leaf_132_clk _01048_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_94_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21727_ _03375_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24446_ clknet_leaf_63_clk net617 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[0\].output_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12460_ _05284_ _05276_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21658_ _03372_ _03386_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12391_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[12\] _05235_
+ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__or2_1
X_20609_ _02378_ _02379_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__and2b_1
X_24377_ clknet_leaf_38_clk _00910_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21589_ _03315_ _03319_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14130_ _06842_ _06844_ VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__nor2_1
X_23328_ net694 _04778_ _04780_ _04769_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14061_ _06648_ _06628_ _06645_ _06626_ VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__nand4_4
XFILLER_0_238_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23259_ net752 _04739_ _04741_ _04730_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13012_ _05793_ _05794_ _05795_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__and3b_1
XTAP_6620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17820_ _10284_ _10288_ _10286_ VGND VGND VPWR VPWR _10327_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_234_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17751_ _10203_ _10217_ _10259_ VGND VGND VPWR VPWR _10260_ sky130_fd_sc_hd__o21a_1
XTAP_5963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14963_ _07626_ VGND VGND VPWR VPWR _07627_ sky130_fd_sc_hd__buf_2
XFILLER_0_55_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_86_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_16
X_16702_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[3\] _08066_ _09262_
+ _09263_ VGND VGND VPWR VPWR _09264_ sky130_fd_sc_hd__a22o_1
XFILLER_0_226_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13914_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _06643_ sky130_fd_sc_hd__clkbuf_4
X_17682_ _10192_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__clkbuf_1
X_14894_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[16\] _07576_ VGND
+ VGND VPWR VPWR _07577_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19421_ _01254_ _01255_ _01228_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_226_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16633_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _09203_ sky130_fd_sc_hd__buf_4
XFILLER_0_202_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13845_ _06567_ _06569_ VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__or2b_1
XFILLER_0_162_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19352_ _01187_ _01188_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[3\]
+ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__a21oi_1
X_16564_ _09137_ _09139_ VGND VGND VPWR VPWR _09140_ sky130_fd_sc_hd__xnor2_1
X_13776_ _06484_ _06480_ _06518_ VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__nand3_1
XFILLER_0_130_1119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18303_ _10768_ _10769_ VGND VGND VPWR VPWR _10770_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15515_ _07619_ _06634_ _08148_ _08142_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__o211a_1
X_12727_ _05535_ _05536_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19283_ _09185_ _11682_ _11685_ _11641_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__o211a_1
X_16495_ _09000_ _09034_ VGND VGND VPWR VPWR _09073_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18234_ _10700_ _10702_ VGND VGND VPWR VPWR _10703_ sky130_fd_sc_hd__xnor2_2
X_15446_ _08086_ _08087_ VGND VGND VPWR VPWR _08088_ sky130_fd_sc_hd__xnor2_2
X_12658_ _05424_ _05469_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18165_ _10635_ _10636_ VGND VGND VPWR VPWR _10637_ sky130_fd_sc_hd__and2_1
X_15377_ _08019_ _08020_ VGND VGND VPWR VPWR _08021_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12589_ _05402_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_clk clknet_4_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17116_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[13\] _09459_ _09417_
+ VGND VGND VPWR VPWR _09667_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14328_ _07035_ _07026_ VGND VGND VPWR VPWR _07037_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18096_ _04858_ VGND VGND VPWR VPWR _10583_ sky130_fd_sc_hd__buf_4
XFILLER_0_29_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold406 _00150_ VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 top_inst.axis_out_inst.out_buff_data\[91\] VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold428 top_inst.axis_out_inst.out_buff_data\[43\] VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold439 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[6\] VGND VGND
+ VPWR VPWR net621 sky130_fd_sc_hd__dlygate4sd3_1
X_17047_ _09597_ _09598_ _09599_ VGND VGND VPWR VPWR _09600_ sky130_fd_sc_hd__nand3_1
XFILLER_0_180_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14259_ _06967_ _06969_ VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_14__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_4_14__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_18998_ _11417_ _11419_ VGND VGND VPWR VPWR _11420_ sky130_fd_sc_hd__nor2_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17949_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[13\] _10367_ VGND
+ VGND VPWR VPWR _10453_ sky130_fd_sc_hd__xnor2_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_77_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_139_1144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20960_ _02727_ _02728_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19619_ _01407_ _01409_ _01408_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_71_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20891_ _02632_ _02659_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__or2_1
XFILLER_0_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22630_ _04288_ _04291_ _04290_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__a21o_1
XFILLER_0_221_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22561_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[17\] _04215_ _04216_
+ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24300_ clknet_leaf_138_clk _00833_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[75\]
+ sky130_fd_sc_hd__dfxtp_1
X_21512_ _03135_ _03208_ _03168_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_173_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22492_ _04161_ _04173_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21443_ _02871_ _02893_ _03140_ _03177_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__a31o_1
X_24231_ clknet_leaf_113_clk _00764_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[16\]\[6\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_17_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24162_ clknet_leaf_13_clk _00695_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_21374_ _02897_ _03062_ _03110_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_47_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23113_ _04655_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__clkbuf_4
X_20325_ _02110_ _02111_ _02109_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24093_ clknet_leaf_99_clk _00626_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23044_ net902 _04616_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__or2_1
X_20256_ _02030_ _02036_ _02046_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_229_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20187_ _10030_ _11687_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__or2_2
XTAP_5226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_68_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_16
XTAP_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23946_ clknet_leaf_90_clk _00479_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_11960_ net783 _04990_ _04991_ _04981_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23877_ clknet_leaf_51_clk _00410_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ net648 _04951_ _04952_ _04942_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13630_ _06195_ _06205_ _06375_ _06376_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_169_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22828_ net499 _09804_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__or2_1
XFILLER_0_211_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13561_ _06305_ _06308_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22759_ _04092_ _04427_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15300_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[10\] _06242_ _07944_
+ _07945_ VGND VGND VPWR VPWR _07946_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12512_ net1026 _05314_ _05329_ _05308_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__o211a_1
X_16280_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[7\] _08862_ VGND
+ VGND VPWR VPWR _08863_ sky130_fd_sc_hd__xnor2_1
X_13492_ _06231_ _06236_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__and2b_1
XFILLER_0_136_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15231_ top_inst.grid_inst.data_path_wires\[6\]\[6\] top_inst.grid_inst.data_path_wires\[6\]\[5\]
+ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _07878_ sky130_fd_sc_hd__and4_1
X_24429_ clknet_leaf_58_clk net719 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].output_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12443_ _05269_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__buf_8
XFILLER_0_168_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15162_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[7\] _07810_ VGND
+ VGND VPWR VPWR _07811_ sky130_fd_sc_hd__xnor2_1
X_12374_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[5\] _05222_
+ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_209_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14113_ _06777_ _06779_ _06826_ VGND VGND VPWR VPWR _06828_ sky130_fd_sc_hd__nand3_1
XFILLER_0_120_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19970_ _01786_ _01787_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__and2_1
X_15093_ _07725_ _07721_ VGND VGND VPWR VPWR _07743_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_240_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14044_ _06723_ _06725_ _06760_ VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__a21oi_1
X_18921_ _11158_ _11140_ _11156_ _11143_ VGND VGND VPWR VPWR _11344_ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18852_ _11275_ _11276_ _11140_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[2\]
+ VGND VGND VPWR VPWR _11277_ sky130_fd_sc_hd__and4bb_1
XTAP_6450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17803_ _10256_ _10254_ VGND VGND VPWR VPWR _10311_ sky130_fd_sc_hd__and2b_1
XTAP_6494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18783_ top_inst.grid_inst.data_path_wires\[13\]\[3\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[13\]\[4\]
+ VGND VGND VPWR VPWR _11210_ sky130_fd_sc_hd__a22o_1
XTAP_5760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15995_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[14\] _08452_ VGND
+ VGND VPWR VPWR _08604_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_59_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_235_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17734_ _10038_ _10047_ _10240_ _10241_ VGND VGND VPWR VPWR _10243_ sky130_fd_sc_hd__nand4_1
XTAP_5793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14946_ _07613_ _07611_ _07614_ _07092_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17665_ _10170_ _10175_ VGND VGND VPWR VPWR _10176_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_221_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14877_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[14\] _07364_ _07280_
+ VGND VGND VPWR VPWR _07561_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16616_ _09188_ VGND VGND VPWR VPWR _09189_ sky130_fd_sc_hd__clkbuf_4
X_19404_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[2\] _11692_ _01238_
+ _01239_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__nand4_4
XFILLER_0_216_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13828_ _06567_ _06569_ VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__xor2_1
X_17596_ _10107_ _10108_ VGND VGND VPWR VPWR _10109_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16547_ _09117_ _09088_ _09122_ VGND VGND VPWR VPWR _09123_ sky130_fd_sc_hd__a21oi_1
X_19335_ _11727_ _11728_ VGND VGND VPWR VPWR _11729_ sky130_fd_sc_hd__nand2_1
X_13759_ _06499_ _06502_ VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19266_ net1018 _11662_ _11675_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16478_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[12\] _08897_ VGND
+ VGND VPWR VPWR _09056_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_922 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18217_ top_inst.grid_inst.data_path_wires\[12\]\[2\] top_inst.grid_inst.data_path_wires\[12\]\[1\]
+ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[4\] VGND VGND VPWR VPWR
+ _10686_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15429_ _07624_ _07824_ _08031_ VGND VGND VPWR VPWR _08071_ sky130_fd_sc_hd__o21a_1
XFILLER_0_170_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19197_ _11610_ _11613_ VGND VGND VPWR VPWR _11614_ sky130_fd_sc_hd__xor2_2
XFILLER_0_182_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18148_ top_inst.grid_inst.data_path_wires\[12\]\[0\] _10600_ _10597_ _10599_ VGND
+ VGND VPWR VPWR _10621_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold203 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[24\] VGND
+ VGND VPWR VPWR net385 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold214 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[0\] VGND VGND
+ VPWR VPWR net396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 _00905_ VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18079_ net928 _10563_ _10576_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__o21a_1
XFILLER_0_229_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold236 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[7\] VGND
+ VGND VPWR VPWR net418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold247 _00038_ VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20110_ _01915_ _01922_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__xnor2_1
Xhold258 top_inst.axis_out_inst.out_buff_data\[10\] VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 top_inst.axis_out_inst.out_buff_data\[122\] VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21090_ _05440_ _02852_ VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__nor2_1
XFILLER_0_229_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20041_ _01855_ _01856_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__nor2_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23800_ clknet_leaf_70_clk _00333_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21992_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _03697_ sky130_fd_sc_hd__buf_2
XFILLER_0_206_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23731_ clknet_leaf_125_clk _00264_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20943_ _02538_ _02539_ _02540_ _02711_ _02709_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__o311a_1
XANTENNA_109 _05313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_240_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23662_ clknet_leaf_132_clk net309 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20874_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[21\] _02470_ VGND
+ VGND VPWR VPWR _02646_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22613_ _04218_ _04289_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__nor2_1
X_23593_ clknet_leaf_101_clk _00126_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22544_ _04200_ _04223_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22475_ top_inst.deskew_buff_inst.col_input\[110\] _05731_ _04156_ _04157_ VGND VGND
+ VPWR VPWR _04158_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24214_ clknet_leaf_17_clk _00747_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_21426_ _03121_ _03152_ _03160_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__a21o_1
XFILLER_0_162_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_241_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24145_ clknet_leaf_18_clk _00678_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_21357_ top_inst.grid_inst.data_path_wires\[17\]\[1\] _02895_ _03052_ VGND VGND VPWR
+ VPWR _03094_ sky130_fd_sc_hd__and3_1
XFILLER_0_241_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20308_ _02070_ _02096_ _05406_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__a21oi_1
X_12090_ net488 _05058_ _05066_ _05062_ VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21288_ _03024_ _03025_ _02992_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__a21oi_1
X_24076_ clknet_leaf_112_clk _00609_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold770 _00976_ VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[17\] VGND VGND
+ VPWR VPWR net963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[13\] VGND VGND
+ VPWR VPWR net974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23027_ net26 _04601_ _04608_ _04606_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__o211a_1
X_20239_ _02027_ _02029_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[1\]
+ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__a21o_1
XFILLER_0_229_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ _07449_ _07454_ _07452_ VGND VGND VPWR VPWR _07486_ sky130_fd_sc_hd__a21o_1
XTAP_5078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[8\] _07866_ VGND
+ VGND VPWR VPWR _08395_ sky130_fd_sc_hd__or2_1
XFILLER_0_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12992_ _05734_ _05759_ _05757_ _05738_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__a22o_1
XTAP_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14731_ _07083_ _07086_ _07417_ _07418_ VGND VGND VPWR VPWR _07419_ sky130_fd_sc_hd__nand4_1
XTAP_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23929_ clknet_leaf_76_clk _00462_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ _04876_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__buf_2
XFILLER_0_197_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _09930_ _09986_ _09968_ VGND VGND VPWR VPWR _09987_ sky130_fd_sc_hd__and3_1
XTAP_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14662_ _07304_ _07275_ VGND VGND VPWR VPWR _07352_ sky130_fd_sc_hd__or2b_1
XTAP_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11874_ _04876_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__buf_2
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _08974_ _08980_ VGND VGND VPWR VPWR _08981_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[7\] _05326_ VGND
+ VGND VPWR VPWR _06361_ sky130_fd_sc_hd__and2_1
XFILLER_0_211_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17381_ _09918_ _09920_ VGND VGND VPWR VPWR _09921_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14593_ _07276_ _07283_ VGND VGND VPWR VPWR _07284_ sky130_fd_sc_hd__xor2_1
XFILLER_0_139_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19120_ _11509_ _11538_ VGND VGND VPWR VPWR _11539_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16332_ _08873_ _08874_ _08913_ VGND VGND VPWR VPWR _08914_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13544_ _06292_ _06277_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19051_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[11\] _11340_ VGND
+ VGND VPWR VPWR _11471_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16263_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[6\] _08809_ _08810_
+ VGND VGND VPWR VPWR _08846_ sky130_fd_sc_hd__a21bo_1
X_13475_ _06226_ _06227_ _05336_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_124_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18002_ _10464_ _10467_ _10503_ VGND VGND VPWR VPWR _10505_ sky130_fd_sc_hd__and3_1
XFILLER_0_164_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15214_ _07821_ _07822_ _07861_ VGND VGND VPWR VPWR _07862_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12426_ net369 _05256_ _05257_ _05247_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__o211a_1
X_16194_ _08770_ _08778_ VGND VGND VPWR VPWR _08779_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_239_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15145_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[6\] _07756_ _07757_
+ VGND VGND VPWR VPWR _07794_ sky130_fd_sc_hd__a21bo_1
X_12357_ net695 _05217_ _05218_ _05208_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_1430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19953_ _01737_ _01745_ _01770_ _01726_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_142_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15076_ _07720_ _07726_ VGND VGND VPWR VPWR _07727_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_227_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12288_ net490 _05178_ _05179_ _05168_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_1097 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14027_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[3\]
+ top_inst.grid_inst.data_path_wires\[3\]\[3\] _06624_ VGND VGND VPWR VPWR _06744_
+ sky130_fd_sc_hd__nand4_2
X_18904_ _11288_ _11327_ VGND VGND VPWR VPWR _11328_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19884_ _01705_ _01702_ _01706_ VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_219_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18835_ _11243_ _11239_ VGND VGND VPWR VPWR _11260_ sky130_fd_sc_hd__or2b_1
XFILLER_0_235_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18766_ _11192_ _11193_ VGND VGND VPWR VPWR _11194_ sky130_fd_sc_hd__nand2_2
X_15978_ _08546_ _08587_ VGND VGND VPWR VPWR _08588_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14929_ _07593_ _07603_ _07594_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17717_ _10224_ _10225_ _05353_ VGND VGND VPWR VPWR _10227_ sky130_fd_sc_hd__a21o_1
XFILLER_0_222_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18697_ top_inst.grid_inst.data_path_wires\[13\]\[4\] VGND VGND VPWR VPWR _11140_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17648_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[5\] _10136_ _10137_
+ VGND VGND VPWR VPWR _10159_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_33_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17579_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[3\] _10091_ _10092_
+ VGND VGND VPWR VPWR _10093_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19318_ _10447_ VGND VGND VPWR VPWR _11714_ sky130_fd_sc_hd__buf_2
X_20590_ _02327_ _02333_ _02364_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19249_ _11655_ _11657_ VGND VGND VPWR VPWR _11663_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22260_ _03947_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21211_ top_inst.grid_inst.data_path_wires\[17\]\[0\] _02891_ _02889_ top_inst.grid_inst.data_path_wires\[17\]\[1\]
+ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22191_ _03841_ _03843_ _03840_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_48_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21142_ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _02891_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21073_ _02821_ _02836_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20024_ _01819_ _01838_ _01839_ _01840_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21975_ _02866_ _02877_ _03685_ _03660_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__o211a_1
Xrebuffer40 net221 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer51 net239 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_240_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer62 net243 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23714_ clknet_leaf_123_clk _00247_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer73 net1119 VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__buf_2
XFILLER_0_16_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20926_ _02503_ _02687_ _02694_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__or3_1
XFILLER_0_194_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23645_ clknet_leaf_123_clk net593 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20857_ _02603_ _02615_ _02628_ VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__nand3_1
XFILLER_0_166_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23576_ clknet_leaf_107_clk _00109_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20788_ _02562_ _02563_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22527_ _04177_ _04207_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_1186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13260_ _06035_ _06036_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__or2_1
X_22458_ _04025_ _04139_ _04140_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__nor3_1
XFILLER_0_33_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12211_ top_inst.axis_out_inst.out_buff_data\[31\] _05129_ VGND VGND VPWR VPWR _05135_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_121_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21409_ _03136_ _03144_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__xnor2_2
X_13191_ top_inst.grid_inst.data_path_wires\[1\]\[2\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__and2b_1
XFILLER_0_150_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22389_ _04071_ _04073_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__xor2_1
XFILLER_0_241_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12142_ net432 _05084_ _05095_ _05088_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__o211a_1
X_24128_ clknet_leaf_117_clk _00661_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_102_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16950_ _09501_ _09504_ VGND VGND VPWR VPWR _09505_ sky130_fd_sc_hd__xor2_1
X_24059_ clknet_leaf_45_clk _00592_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_21_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12073_ net514 _05045_ _05056_ _05049_ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__o211a_1
X_15901_ _08469_ _08471_ _08467_ VGND VGND VPWR VPWR _08513_ sky130_fd_sc_hd__a21oi_1
X_16881_ _09375_ _09383_ _09382_ VGND VGND VPWR VPWR _09438_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15832_ _08149_ _08164_ _08161_ top_inst.grid_inst.data_path_wires\[7\]\[7\] VGND
+ VGND VPWR VPWR _08445_ sky130_fd_sc_hd__a22o_1
X_18620_ _10969_ _11078_ VGND VGND VPWR VPWR _11079_ sky130_fd_sc_hd__nor2_1
XFILLER_0_205_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _08376_ _08377_ VGND VGND VPWR VPWR _08378_ sky130_fd_sc_hd__nor2_1
X_18551_ _10979_ _10980_ _10982_ VGND VGND VPWR VPWR _11012_ sky130_fd_sc_hd__or3_1
XFILLER_0_235_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12975_ _05765_ _05294_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__or2_1
XTAP_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_234_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14714_ _06848_ _07401_ _07402_ _07092_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__o211a_1
X_17502_ _10029_ _07611_ _10031_ _10024_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__o211a_1
XTAP_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ net558 _04964_ _04972_ _04968_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__o211a_1
X_18482_ _10942_ _10944_ VGND VGND VPWR VPWR _10945_ sky130_fd_sc_hd__xor2_1
XFILLER_0_197_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15694_ _08276_ _08281_ VGND VGND VPWR VPWR _08310_ sky130_fd_sc_hd__nor2_1
XTAP_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17433_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[27\] _05316_ VGND
+ VGND VPWR VPWR _09971_ sky130_fd_sc_hd__or2_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[7\] _07290_ _07073_
+ _07087_ VGND VGND VPWR VPWR _07335_ sky130_fd_sc_hd__a22o_1
XFILLER_0_184_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ net860 _04925_ _04933_ _04929_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__o211a_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17364_ _09880_ _09904_ VGND VGND VPWR VPWR _09905_ sky130_fd_sc_hd__xnor2_2
X_14576_ _07221_ _07223_ _07219_ VGND VGND VPWR VPWR _07268_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_172_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11788_ top_inst.axis_out_inst.out_buff_data\[73\] _04890_ VGND VGND VPWR VPWR _04894_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_83_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16315_ _08894_ _08896_ VGND VGND VPWR VPWR _08897_ sky130_fd_sc_hd__nor2_4
X_19103_ _11164_ _11145_ _11521_ VGND VGND VPWR VPWR _11522_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13527_ _06271_ _06276_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__xnor2_2
X_17295_ _09834_ _09838_ VGND VGND VPWR VPWR _09839_ sky130_fd_sc_hd__xor2_2
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19034_ _11453_ _11454_ VGND VGND VPWR VPWR _11455_ sky130_fd_sc_hd__xnor2_1
X_16246_ _08197_ _08829_ VGND VGND VPWR VPWR _08830_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13458_ _06214_ _05773_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12409_ _05142_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_113_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16177_ _08738_ _08758_ VGND VGND VPWR VPWR _08762_ sky130_fd_sc_hd__nor2_1
X_13389_ _06159_ _06160_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__nand2_1
Xoutput105 net105 VGND VGND VPWR VPWR output_tdata[45] sky130_fd_sc_hd__buf_2
XFILLER_0_23_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput116 net116 VGND VGND VPWR VPWR output_tdata[55] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput127 net127 VGND VGND VPWR VPWR output_tdata[65] sky130_fd_sc_hd__clkbuf_4
Xoutput138 net138 VGND VGND VPWR VPWR output_tdata[75] sky130_fd_sc_hd__clkbuf_4
X_15128_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[6\] _07777_ _06701_
+ VGND VGND VPWR VPWR _07778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput149 net149 VGND VGND VPWR VPWR output_tdata[85] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19936_ _01755_ _01756_ _06682_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__a21o_1
X_15059_ _07695_ _07699_ VGND VGND VPWR VPWR _07710_ sky130_fd_sc_hd__and2b_1
XFILLER_0_120_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19867_ _01679_ _01680_ _01690_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_128_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_235_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18818_ _11239_ _11243_ VGND VGND VPWR VPWR _11244_ sky130_fd_sc_hd__xnor2_2
X_19798_ _11722_ _01624_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18749_ _11154_ _11130_ VGND VGND VPWR VPWR _11178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21760_ _03460_ _03483_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__or2_1
XFILLER_0_176_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20711_ _02135_ _02489_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__and2_1
XFILLER_0_187_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21691_ _03402_ _03417_ _03418_ _05309_ _04861_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_86_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23430_ net290 _04827_ _04836_ _04831_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20642_ _02390_ _02418_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23361_ net44 _04792_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__or2_1
X_20573_ _02318_ _02320_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22312_ _03982_ _03998_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23292_ net138 _04753_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22243_ _03887_ _03926_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22174_ _03690_ _03703_ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21125_ _02878_ _02869_ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21056_ _02794_ _02796_ _02820_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_195_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20007_ _01652_ _01751_ _01793_ _01820_ _01823_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__a41o_4
XFILLER_0_195_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_241_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12760_ _05565_ _05568_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__nand2_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21958_ _02885_ _02883_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20909_ _02678_ _02679_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__or2_1
X_12691_ _05496_ _05501_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21889_ top_inst.deskew_buff_inst.col_input\[90\] _05325_ VGND VGND VPWR VPWR _03608_
+ sky130_fd_sc_hd__and2_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _07074_ _07061_ _07065_ _07070_ VGND VGND VPWR VPWR _07126_ sky130_fd_sc_hd__a22o_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23628_ clknet_leaf_102_clk net275 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_204_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14361_ _07066_ _06641_ VGND VGND VPWR VPWR _07067_ sky130_fd_sc_hd__or2_1
XFILLER_0_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_944 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23559_ clknet_leaf_100_clk net806 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16100_ _08693_ _08684_ VGND VGND VPWR VPWR _08694_ sky130_fd_sc_hd__or2_1
Xinput18 input_tdata[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_4
XFILLER_0_108_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13312_ _06083_ _06084_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__nor2_1
Xinput29 input_tdata[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_4
X_17080_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[13\] _09631_ VGND
+ VGND VPWR VPWR _09632_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14292_ _06965_ _06969_ _07001_ VGND VGND VPWR VPWR _07002_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16031_ _08612_ _08613_ _08610_ VGND VGND VPWR VPWR _08639_ sky130_fd_sc_hd__o21a_1
XFILLER_0_243_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13243_ _06015_ _06019_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_1015 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13174_ _05943_ _05952_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_209_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12125_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[26\] _05076_
+ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17982_ _10450_ _10449_ VGND VGND VPWR VPWR _10485_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19721_ _01522_ _01548_ _01549_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__and3_1
X_16933_ _09487_ _09488_ VGND VGND VPWR VPWR _09489_ sky130_fd_sc_hd__and2_1
X_12056_ net266 _05036_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__or2_1
XFILLER_0_237_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19652_ _01479_ _01481_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__xnor2_1
X_16864_ _09415_ _09420_ VGND VGND VPWR VPWR _09421_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_244_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_204_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18603_ _11061_ _11043_ VGND VGND VPWR VPWR _11063_ sky130_fd_sc_hd__or2b_1
X_15815_ _08426_ _08428_ VGND VGND VPWR VPWR _08429_ sky130_fd_sc_hd__nor2_1
X_16795_ _09352_ _09353_ VGND VGND VPWR VPWR _09354_ sky130_fd_sc_hd__and2_1
X_19583_ _01406_ _01413_ _01414_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__nand3_2
XFILLER_0_204_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15746_ _08163_ _08164_ _08161_ _08147_ VGND VGND VPWR VPWR _08361_ sky130_fd_sc_hd__a22o_1
X_18534_ _10961_ _10962_ _10994_ VGND VGND VPWR VPWR _10996_ sky130_fd_sc_hd__and3_1
X_12958_ _05736_ _05306_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11909_ net561 _04951_ _04962_ _04955_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__o211a_1
X_18465_ _10926_ _10925_ VGND VGND VPWR VPWR _10928_ sky130_fd_sc_hd__and2b_1
X_15677_ _08283_ _08292_ VGND VGND VPWR VPWR _08294_ sky130_fd_sc_hd__or2_1
X_12889_ _05664_ _05667_ _05693_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__o21ai_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14628_ _07276_ _07283_ _07317_ VGND VGND VPWR VPWR _07318_ sky130_fd_sc_hd__a21bo_2
X_17416_ _09624_ _09953_ VGND VGND VPWR VPWR _09954_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18396_ _10585_ _10610_ _10804_ _10803_ VGND VGND VPWR VPWR _10861_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17347_ _09850_ _09887_ VGND VGND VPWR VPWR _09888_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14559_ _07235_ _07249_ _07250_ VGND VGND VPWR VPWR _07251_ sky130_fd_sc_hd__nand3_1
XFILLER_0_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17278_ _09782_ _09801_ VGND VGND VPWR VPWR _09823_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16229_ _08808_ _08812_ VGND VGND VPWR VPWR _08813_ sky130_fd_sc_hd__xor2_1
X_19017_ top_inst.grid_inst.data_path_wires\[13\]\[7\] _11158_ _11156_ VGND VGND VPWR
+ VPWR _11438_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19919_ _01561_ _01739_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22930_ net994 _04548_ _04552_ _04551_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22861_ net828 _04504_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__or2_1
XFILLER_0_211_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24600_ clknet_leaf_24_clk _01133_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_39_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21812_ _03515_ _03533_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_223_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22792_ _04408_ _04458_ _04460_ _04440_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24531_ clknet_leaf_129_clk _01064_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dfxtp_4
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21743_ _03438_ _03440_ _03463_ _03467_ _03462_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__a32oi_4
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24462_ clknet_leaf_57_clk _00995_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21674_ _03394_ _03399_ _03392_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__o21a_1
XFILLER_0_163_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23413_ net1014 _04588_ _04826_ _04819_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20625_ _02003_ _02018_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__nand2_2
X_24393_ clknet_leaf_38_clk net853 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23344_ net163 _04779_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20556_ _02297_ _02299_ _02337_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__nand3_1
XFILLER_0_225_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23275_ net130 _04740_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__or2_1
X_20487_ _02228_ _02232_ net178 _02270_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__o31ai_2
X_22226_ _03897_ _03914_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_225_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22157_ _03812_ _03819_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__or2b_1
XFILLER_0_160_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21108_ _02866_ _11133_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__or2_1
X_22088_ _03686_ _03703_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13930_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[7\] _06641_ VGND
+ VGND VPWR VPWR _06654_ sky130_fd_sc_hd__or2_1
X_21039_ net997 _02491_ _02802_ _02804_ _01863_ VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__o221a_1
XFILLER_0_156_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13861_ _06600_ _06601_ VGND VGND VPWR VPWR _06602_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15600_ top_inst.grid_inst.data_path_wires\[7\]\[3\] top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[1\]
+ _08154_ top_inst.grid_inst.data_path_wires\[7\]\[4\] VGND VGND VPWR VPWR _08219_
+ sky130_fd_sc_hd__a22o_1
X_12812_ _05614_ _05618_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__nor2_1
XFILLER_0_236_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16580_ _09152_ _09154_ VGND VGND VPWR VPWR _09155_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_201_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13792_ _06523_ _06498_ _06534_ VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__a21o_1
XFILLER_0_232_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15531_ _08159_ _07641_ VGND VGND VPWR VPWR _08160_ sky130_fd_sc_hd__or2_1
X_12743_ _05550_ _05551_ _05525_ _05526_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__o211a_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ top_inst.grid_inst.data_path_wires\[12\]\[5\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[0\] _10591_ VGND VGND
+ VPWR VPWR _10718_ sky130_fd_sc_hd__a22o_1
X_15462_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[14\] _07924_ _07844_
+ VGND VGND VPWR VPWR _08103_ sky130_fd_sc_hd__a21o_1
X_12674_ _05424_ _05469_ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__nand2_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _09727_ _09737_ VGND VGND VPWR VPWR _09749_ sky130_fd_sc_hd__or2_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _07070_ _07061_ _07109_ VGND VGND VPWR VPWR _07110_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18181_ _10650_ _10651_ VGND VGND VPWR VPWR _10652_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15393_ _07990_ _07993_ _07992_ VGND VGND VPWR VPWR _08036_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_5_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17132_ _09681_ _09682_ VGND VGND VPWR VPWR _09683_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14344_ _06995_ _07038_ _07036_ VGND VGND VPWR VPWR _07052_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17063_ _09584_ _09615_ VGND VGND VPWR VPWR _09616_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14275_ _06907_ _06952_ _06950_ VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16014_ _08620_ _08621_ _08265_ VGND VGND VPWR VPWR _08623_ sky130_fd_sc_hd__o21a_1
X_13226_ _06002_ _06003_ _05328_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__a21o_1
XFILLER_0_243_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13157_ top_inst.grid_inst.data_path_wires\[1\]\[5\] _05746_ _05765_ _05763_ VGND
+ VGND VPWR VPWR _05936_ sky130_fd_sc_hd__nand4_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12108_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[18\] _05076_
+ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__or2_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _05864_ _05867_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__nor2_1
X_17965_ _10467_ _10468_ VGND VGND VPWR VPWR _10469_ sky130_fd_sc_hd__nand2_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19704_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[5\] _11707_ VGND
+ VGND VPWR VPWR _01533_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16916_ _09361_ net223 _09201_ _09213_ VGND VGND VPWR VPWR _09472_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12039_ net861 _05031_ _05037_ _05035_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17896_ _10357_ _10360_ _10400_ _07439_ VGND VGND VPWR VPWR _10402_ sky130_fd_sc_hd__a31o_1
XFILLER_0_217_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19635_ _01464_ _01465_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__or2_4
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16847_ _09403_ _09404_ VGND VGND VPWR VPWR _09405_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19566_ _11688_ _11705_ _01361_ _01360_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__a31o_1
X_16778_ _09213_ _09186_ _09192_ _09211_ VGND VGND VPWR VPWR _09337_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_220_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18517_ _10975_ _10977_ _10978_ VGND VGND VPWR VPWR _10979_ sky130_fd_sc_hd__nor3_1
XFILLER_0_158_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_1082 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15729_ _08342_ _08343_ _06404_ VGND VGND VPWR VPWR _08345_ sky130_fd_sc_hd__a21o_1
X_19497_ _01328_ _01329_ net198 _01268_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18448_ _10882_ _10883_ _10910_ VGND VGND VPWR VPWR _10912_ sky130_fd_sc_hd__nand3_1
XFILLER_0_185_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18379_ _10798_ _10800_ _10842_ VGND VGND VPWR VPWR _10844_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20410_ _02149_ _02150_ _02151_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_209_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21390_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[9\] _03080_ VGND
+ VGND VPWR VPWR _03126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20341_ _02093_ _02092_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23060_ net10 _04615_ _04626_ _04619_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__o211a_1
X_20272_ _02041_ _02059_ _02060_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__and3_1
XFILLER_0_222_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22011_ _03690_ _05270_ _03710_ _03702_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__o211a_1
XTAP_6109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23962_ clknet_leaf_89_clk _00495_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_192_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22913_ top_inst.skew_buff_inst.row\[2\].output_reg\[4\] _04530_ VGND VGND VPWR VPWR
+ _04542_ sky130_fd_sc_hd__or2_1
XFILLER_0_230_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23893_ clknet_leaf_52_clk _00426_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22844_ top_inst.skew_buff_inst.row\[3\].output_reg\[6\] _03691_ VGND VGND VPWR VPWR
+ _04503_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_233_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22775_ _04410_ _04430_ _04428_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24514_ clknet_leaf_132_clk _01047_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_109_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21726_ _03447_ _03451_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_164_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24445_ clknet_leaf_63_clk net1020 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[0\].output_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21657_ _03384_ _03385_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_1408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20608_ _02385_ _02388_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__nand2_1
X_24376_ clknet_leaf_39_clk net851 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].output_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12390_ net535 _05230_ _05237_ _05234_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21588_ _03317_ _03318_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23327_ net155 _04779_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__or2_1
X_20539_ _02316_ _02321_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14060_ top_inst.grid_inst.data_path_wires\[3\]\[4\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[3\]
+ _06626_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _06776_ sky130_fd_sc_hd__a22o_1
X_23258_ net122 _04740_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__or2_1
XFILLER_0_240_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13011_ _05777_ _05781_ _05792_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__or3_1
X_22209_ _03707_ _03688_ _03705_ _03690_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23189_ net89 _04701_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__or2_1
XTAP_6621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14962_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _07626_ sky130_fd_sc_hd__buf_2
X_17750_ _10204_ _10216_ VGND VGND VPWR VPWR _10259_ sky130_fd_sc_hd__nand2_1
XFILLER_0_233_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16701_ _09243_ _09261_ _05399_ VGND VGND VPWR VPWR _09263_ sky130_fd_sc_hd__a21oi_1
XTAP_5997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13913_ _06622_ _06204_ _06642_ _06639_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14893_ _05731_ VGND VGND VPWR VPWR _07576_ sky130_fd_sc_hd__buf_8
X_17681_ _09661_ _10191_ VGND VGND VPWR VPWR _10192_ sky130_fd_sc_hd__and2_1
XFILLER_0_226_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_242_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19420_ _01228_ _01254_ _01255_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__and3_1
X_16632_ _09201_ VGND VGND VPWR VPWR _09202_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13844_ _06585_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19351_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[3\] _01187_ _01188_
+ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__and3_1
X_16563_ _09101_ _09102_ _09138_ VGND VGND VPWR VPWR _09139_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13775_ _06484_ _06480_ _06518_ VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__a21o_1
XFILLER_0_202_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18302_ top_inst.grid_inst.data_path_wires\[12\]\[0\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _10769_ sky130_fd_sc_hd__and2b_1
X_12726_ _05293_ _05288_ _05297_ _05301_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__and4_1
X_15514_ _08147_ _08140_ VGND VGND VPWR VPWR _08148_ sky130_fd_sc_hd__or2_1
X_16494_ _09032_ _09071_ VGND VGND VPWR VPWR _09072_ sky130_fd_sc_hd__xor2_2
X_19282_ _11684_ _11150_ VGND VGND VPWR VPWR _11685_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15445_ _08043_ _08047_ _08045_ VGND VGND VPWR VPWR _08087_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_66_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18233_ _10668_ _10669_ _10701_ VGND VGND VPWR VPWR _10702_ sky130_fd_sc_hd__a21o_1
X_12657_ _05462_ _05468_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15376_ _08016_ _08018_ VGND VGND VPWR VPWR _08020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18164_ _10628_ _10634_ VGND VGND VPWR VPWR _10636_ sky130_fd_sc_hd__nand2_1
X_12588_ _05352_ _05401_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17115_ _09627_ _09652_ _09650_ VGND VGND VPWR VPWR _09666_ sky130_fd_sc_hd__a21o_1
X_14327_ _07026_ _07035_ VGND VGND VPWR VPWR _07036_ sky130_fd_sc_hd__and2b_1
XFILLER_0_170_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18095_ _10027_ _08663_ _10582_ _10448_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold407 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[0\] VGND
+ VGND VPWR VPWR net589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold418 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[4\] VGND
+ VGND VPWR VPWR net600 sky130_fd_sc_hd__dlygate4sd3_1
X_17046_ _09361_ _09210_ net203 _09213_ VGND VGND VPWR VPWR _09599_ sky130_fd_sc_hd__a2bb2o_1
X_14258_ _06635_ _06650_ _06968_ VGND VGND VPWR VPWR _06969_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold429 top_inst.deskew_buff_inst.col_input\[78\] VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13209_ _05748_ _05746_ _05765_ _05763_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14189_ _06897_ _06901_ VGND VGND VPWR VPWR _06902_ sky130_fd_sc_hd__xnor2_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _11335_ _11365_ _11418_ VGND VGND VPWR VPWR _11419_ sky130_fd_sc_hd__a21oi_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[12\] _10367_ _10283_
+ VGND VGND VPWR VPWR _10452_ sky130_fd_sc_hd__a21o_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17879_ _10339_ _10341_ _10340_ VGND VGND VPWR VPWR _10385_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_75_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19618_ _01446_ _01447_ _01445_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20890_ _01819_ _02660_ _02661_ _02035_ VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19549_ _01346_ _01381_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_959 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22560_ _04217_ _04221_ _04220_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21511_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[11\] _03122_ _03123_
+ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__a21o_1
X_22491_ _04170_ _04172_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_228_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24230_ clknet_leaf_113_clk _00763_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[16\]\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_133_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21442_ top_inst.grid_inst.data_path_wires\[17\]\[3\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[6\]
+ _03138_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24161_ clknet_leaf_13_clk _00694_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21373_ _03061_ _03060_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__and2b_1
XFILLER_0_114_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23112_ _04654_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20324_ _02109_ _02110_ _02111_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__nand3_1
X_24092_ clknet_leaf_99_clk _00625_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold930 top_inst.axis_in_inst.inbuf_bus\[7\] VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23043_ net2 _04615_ _04617_ _04606_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__o211a_1
X_20255_ _02044_ _02045_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__and2b_1
XFILLER_0_229_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20186_ _01992_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__buf_4
XTAP_5216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23945_ clknet_leaf_85_clk _00478_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23876_ clknet_leaf_62_clk _00409_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11890_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[21\] _04943_
+ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__or2_1
XFILLER_0_233_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22827_ _04487_ _04492_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_233_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13560_ _06305_ _06308_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__and2_1
X_22758_ _04218_ _04427_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12511_ _05320_ _05322_ _05328_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__a21o_1
XFILLER_0_183_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21709_ _03414_ _03435_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__nand2_1
X_13491_ _05353_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_125_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22689_ _04334_ _04338_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15230_ _07619_ _07635_ _07633_ _07621_ VGND VGND VPWR VPWR _07877_ sky130_fd_sc_hd__a22o_1
X_24428_ clknet_leaf_54_clk net703 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].output_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12442_ _05268_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__buf_6
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15161_ _07808_ _07809_ VGND VGND VPWR VPWR _07810_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24359_ clknet_leaf_30_clk _00892_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[118\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12373_ net912 _05217_ _05227_ _05221_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__o211a_1
X_14112_ _06777_ _06779_ _06826_ VGND VGND VPWR VPWR _06827_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15092_ _07729_ _07731_ VGND VGND VPWR VPWR _07742_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_239_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14043_ _06707_ _06722_ VGND VGND VPWR VPWR _06760_ sky130_fd_sc_hd__nor2_1
X_18920_ _11336_ _11342_ VGND VGND VPWR VPWR _11343_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18851_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[3\]
+ top_inst.grid_inst.data_path_wires\[13\]\[3\] top_inst.grid_inst.data_path_wires\[13\]\[2\]
+ VGND VGND VPWR VPWR _11276_ sky130_fd_sc_hd__and4_1
XFILLER_0_101_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17802_ _10289_ _10309_ VGND VGND VPWR VPWR _10310_ sky130_fd_sc_hd__xnor2_1
XTAP_6473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18782_ _11209_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__clkbuf_1
XTAP_6495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15994_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[13\] _08452_ _08373_
+ VGND VGND VPWR VPWR _08603_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17733_ _10038_ _10047_ _10240_ _10241_ VGND VGND VPWR VPWR _10242_ sky130_fd_sc_hd__a22o_1
X_14945_ _04865_ _07333_ VGND VGND VPWR VPWR _07614_ sky130_fd_sc_hd__nand2_1
XFILLER_0_234_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17664_ _10173_ _10174_ VGND VGND VPWR VPWR _10175_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14876_ _07526_ _07537_ VGND VGND VPWR VPWR _07560_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_216_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19403_ _11697_ _11693_ net190 _11687_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__nand4_4
XFILLER_0_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16615_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _09188_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13827_ _06496_ _06533_ _06568_ VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_159_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17595_ _10032_ _10029_ _10044_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _10108_ sky130_fd_sc_hd__nand4_1
XFILLER_0_216_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19334_ _11725_ _11726_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[2\]
+ VGND VGND VPWR VPWR _11728_ sky130_fd_sc_hd__a21o_1
X_16546_ _09007_ _09121_ VGND VGND VPWR VPWR _09122_ sky130_fd_sc_hd__xor2_1
X_13758_ _06500_ _06461_ _06501_ VGND VGND VPWR VPWR _06502_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12709_ _05472_ _05474_ _05518_ _05519_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_45_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19265_ net960 _11662_ _11675_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16477_ _08932_ _09005_ _08967_ VGND VGND VPWR VPWR _09055_ sky130_fd_sc_hd__o21ba_2
X_13689_ _06383_ _06392_ _06434_ VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18216_ _10585_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[2\] VGND
+ VGND VPWR VPWR _10685_ sky130_fd_sc_hd__nand2_1
XFILLER_0_171_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15428_ _07990_ _08032_ _08033_ VGND VGND VPWR VPWR _08070_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19196_ _11572_ _11611_ _11612_ VGND VGND VPWR VPWR _11613_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_72_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15359_ _08001_ _08002_ VGND VGND VPWR VPWR _08003_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18147_ net996 _10616_ _10619_ _10620_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold204 _00159_ VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _00934_ VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18078_ net956 _10563_ _10576_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__o21a_1
Xhold226 top_inst.deskew_buff_inst.col_input\[2\] VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold237 _00174_ VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold248 top_inst.deskew_buff_inst.col_input\[90\] VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17029_ _09581_ _09540_ _09575_ VGND VGND VPWR VPWR _09582_ sky130_fd_sc_hd__a21o_1
Xhold259 top_inst.deskew_buff_inst.col_input\[120\] VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20040_ _01827_ _01832_ _01851_ _01806_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21991_ _02878_ _02877_ _03696_ _03660_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23730_ clknet_leaf_125_clk net496 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20942_ _02570_ _02633_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__nor2_1
XFILLER_0_178_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23661_ clknet_leaf_135_clk _00194_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20873_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[21\] _02468_ VGND
+ VGND VPWR VPWR _02645_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22612_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[20\] _04163_ VGND
+ VGND VPWR VPWR _04289_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23592_ clknet_leaf_101_clk _00125_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22543_ _04217_ _04222_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__xor2_2
XFILLER_0_9_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22474_ _04152_ _04155_ _05311_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24213_ clknet_leaf_118_clk _00746_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_21425_ _03149_ _03151_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_241_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24144_ clknet_leaf_18_clk _00677_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_60_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21356_ _03089_ _03092_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20307_ _02094_ _02095_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_198_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24075_ clknet_leaf_114_clk _00608_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold760 top_inst.axis_in_inst.inbuf_bus\[25\] VGND VGND VPWR VPWR net942 sky130_fd_sc_hd__dlygate4sd3_1
X_21287_ _02992_ _03024_ _03025_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__and3_1
Xhold771 top_inst.deskew_buff_inst.col_input\[89\] VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__buf_1
Xhold782 top_inst.deskew_buff_inst.col_input\[105\] VGND VGND VPWR VPWR net964 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_130_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23026_ net979 _04603_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold793 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[23\] VGND VGND
+ VPWR VPWR net975 sky130_fd_sc_hd__dlygate4sd3_1
X_20238_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[1\] _02027_ _02029_
+ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__nand3_2
XTAP_5002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20169_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[31\] _01976_ VGND
+ VGND VPWR VPWR _01979_ sky130_fd_sc_hd__xnor2_1
XTAP_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _05738_ _05759_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__nand2_1
XTAP_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_1075 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14730_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[7\] _07378_ _07082_
+ _07087_ VGND VGND VPWR VPWR _07418_ sky130_fd_sc_hd__a22o_1
XTAP_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11942_ net1012 _04977_ _04980_ _04981_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23928_ clknet_leaf_76_clk _00461_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _07302_ _07303_ VGND VGND VPWR VPWR _07351_ sky130_fd_sc_hd__or2b_1
XFILLER_0_135_1351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23859_ clknet_leaf_77_clk _00392_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_54_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11873_ net818 _04938_ _04941_ _04942_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__o211a_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16400_ _08976_ _08979_ VGND VGND VPWR VPWR _08980_ sky130_fd_sc_hd__xor2_1
XFILLER_0_156_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ _06320_ _06322_ _06358_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__o21ai_2
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _07277_ _07282_ VGND VGND VPWR VPWR _07283_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17380_ _09919_ _09899_ VGND VGND VPWR VPWR _09920_ sky130_fd_sc_hd__nor2_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16331_ _08910_ _08912_ VGND VGND VPWR VPWR _08913_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13543_ _06270_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__inv_2
XFILLER_0_211_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16262_ _08832_ _08844_ VGND VGND VPWR VPWR _08845_ sky130_fd_sc_hd__xnor2_1
X_19050_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[10\] _11469_ _11387_
+ VGND VGND VPWR VPWR _11470_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13474_ _06181_ _06205_ _06225_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__and3_1
XFILLER_0_164_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15213_ _07858_ _07860_ VGND VGND VPWR VPWR _07861_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18001_ _10464_ _10467_ _10503_ VGND VGND VPWR VPWR _10504_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12425_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[27\] _05248_
+ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16193_ _08771_ _08777_ VGND VGND VPWR VPWR _08778_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_164_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15144_ _07780_ _07792_ VGND VGND VPWR VPWR _07793_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12356_ net304 _05209_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19952_ _01760_ _01771_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__xnor2_2
X_15075_ _07721_ _07725_ VGND VGND VPWR VPWR _07726_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12287_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[31\] _05169_
+ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__or2_1
XFILLER_0_239_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14026_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[3\]\[3\]
+ top_inst.grid_inst.data_path_wires\[3\]\[2\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[4\]
+ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__a22o_1
X_18903_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[7\] _11326_ VGND
+ VGND VPWR VPWR _11327_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_226_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19883_ _01689_ _01681_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__or2b_1
XFILLER_0_219_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18834_ _11247_ _11249_ VGND VGND VPWR VPWR _11259_ sky130_fd_sc_hd__nand2_1
XTAP_6270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18765_ _11156_ _11154_ _11132_ _11130_ VGND VGND VPWR VPWR _11193_ sky130_fd_sc_hd__nand4_4
XFILLER_0_101_1085 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15977_ _08585_ _08586_ VGND VGND VPWR VPWR _08587_ sky130_fd_sc_hd__and2_1
XTAP_5591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17716_ _10224_ _10225_ VGND VGND VPWR VPWR _10226_ sky130_fd_sc_hd__nor2_1
X_14928_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[25\] _07576_ VGND
+ VGND VPWR VPWR _07603_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18696_ _10585_ _10584_ _11139_ _11137_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__o211a_1
XTAP_4890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17647_ _10133_ _10141_ VGND VGND VPWR VPWR _10158_ sky130_fd_sc_hd__and2_1
X_14859_ _07542_ _07543_ VGND VGND VPWR VPWR _07544_ sky130_fd_sc_hd__or2b_1
XFILLER_0_203_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17578_ _10029_ _10027_ _10044_ _10042_ VGND VGND VPWR VPWR _10092_ sky130_fd_sc_hd__nand4_1
XFILLER_0_147_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19317_ _11711_ _11712_ _08181_ VGND VGND VPWR VPWR _11713_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_129_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16529_ _09063_ _09065_ VGND VGND VPWR VPWR _09106_ sky130_fd_sc_hd__or2b_1
XFILLER_0_85_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19248_ _05313_ VGND VGND VPWR VPWR _11662_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19179_ _11594_ _11595_ VGND VGND VPWR VPWR _11596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21210_ _02866_ _02887_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_223_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22190_ _03838_ _03879_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21141_ _02868_ _02881_ _02890_ _02880_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21072_ _02834_ _02835_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20023_ _10447_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21974_ _03684_ _02869_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__or2_1
XFILLER_0_240_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer30 net211 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer41 _09196_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23713_ clknet_leaf_123_clk _00246_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_234_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer52 net239 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20925_ _02503_ _02687_ _02694_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__o21ai_1
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer63 net243 VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__clkbuf_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer74 _09559_ VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__clkbuf_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23644_ clknet_leaf_126_clk net358 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20856_ _02603_ _02615_ _02628_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23575_ clknet_leaf_104_clk _00108_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_20787_ _02527_ _02547_ _02561_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__nand3_1
XFILLER_0_64_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22526_ _04205_ _04206_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22457_ _03695_ _03711_ _03709_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12210_ net339 _05123_ _05134_ _05128_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__o211a_1
X_21408_ _03141_ _03143_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__xor2_2
X_13190_ _05967_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22388_ _03693_ _03709_ _04029_ _04072_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12141_ top_inst.axis_out_inst.out_buff_data\[1\] _05089_ VGND VGND VPWR VPWR _05095_
+ sky130_fd_sc_hd__or2_1
X_24127_ clknet_leaf_118_clk _00660_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21339_ _03045_ _03048_ _03046_ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_202_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_241_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24058_ clknet_leaf_83_clk _00591_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_12072_ net478 _05050_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__or2_1
Xhold590 top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[2\] VGND VGND
+ VPWR VPWR net772 sky130_fd_sc_hd__dlygate4sd3_1
X_23009_ top_inst.skew_buff_inst.row\[0\].output_reg\[5\] _04596_ VGND VGND VPWR VPWR
+ _04597_ sky130_fd_sc_hd__or2_1
X_15900_ _08477_ _08511_ VGND VGND VPWR VPWR _08512_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_194_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16880_ _09434_ _09435_ _09427_ VGND VGND VPWR VPWR _09437_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15831_ top_inst.grid_inst.data_path_wires\[7\]\[7\] _08164_ _08161_ VGND VGND VPWR
+ VPWR _08444_ sky130_fd_sc_hd__and3_1
XFILLER_0_244_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_232_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18550_ _11006_ _11010_ VGND VGND VPWR VPWR _11011_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_232_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12974_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _05765_ sky130_fd_sc_hd__clkbuf_4
XTAP_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15762_ _08318_ _08320_ _08375_ VGND VGND VPWR VPWR _08377_ sky130_fd_sc_hd__and3_1
XTAP_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17501_ _10030_ _09202_ VGND VGND VPWR VPWR _10031_ sky130_fd_sc_hd__or2_1
XTAP_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_971 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14713_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[10\] _06168_ VGND
+ VGND VPWR VPWR _07402_ sky130_fd_sc_hd__or2_1
XTAP_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ net378 _04969_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__or2_1
X_18481_ _10895_ _10902_ _10943_ VGND VGND VPWR VPWR _10944_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_234_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _08309_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17432_ _09932_ _09946_ _09968_ VGND VGND VPWR VPWR _09970_ sky130_fd_sc_hd__and3_1
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14644_ _07241_ _07242_ _07069_ _07333_ VGND VGND VPWR VPWR _07334_ sky130_fd_sc_hd__or4_4
X_11856_ net360 _04930_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__or2_1
XFILLER_0_234_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14575_ _07265_ _07266_ VGND VGND VPWR VPWR _07267_ sky130_fd_sc_hd__nor2_1
X_17363_ _09902_ _09903_ VGND VGND VPWR VPWR _09904_ sky130_fd_sc_hd__xor2_2
XFILLER_0_28_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11787_ net803 _04885_ _04893_ _04889_ VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19102_ _11351_ _11143_ VGND VGND VPWR VPWR _11521_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16314_ _08895_ VGND VGND VPWR VPWR _08896_ sky130_fd_sc_hd__buf_4
XFILLER_0_83_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13526_ _06272_ _06275_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__xor2_2
X_17294_ _09836_ _09837_ VGND VGND VPWR VPWR _09838_ sky130_fd_sc_hd__and2_2
XFILLER_0_32_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19033_ _11393_ _11412_ _11410_ VGND VGND VPWR VPWR _11454_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16245_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[6\] _08828_ _08307_
+ VGND VGND VPWR VPWR _08829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13457_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _06214_ sky130_fd_sc_hd__buf_2
XFILLER_0_88_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12408_ net329 _05243_ _05246_ _05247_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__o211a_1
XFILLER_0_242_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16176_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[4\] _07048_ _08760_
+ _08761_ _07708_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__o221a_1
X_13388_ _06159_ _06160_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__or2_1
Xoutput106 net106 VGND VGND VPWR VPWR output_tdata[46] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_224_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput117 net117 VGND VGND VPWR VPWR output_tdata[56] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput128 net128 VGND VGND VPWR VPWR output_tdata[66] sky130_fd_sc_hd__clkbuf_4
X_15127_ _07775_ _07776_ VGND VGND VPWR VPWR _07777_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12339_ net540 _05204_ _05207_ _05208_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__o211a_1
Xoutput139 net139 VGND VGND VPWR VPWR output_tdata[76] sky130_fd_sc_hd__clkbuf_4
X_19935_ _01749_ _01754_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__or2_1
X_15058_ _07684_ _07703_ VGND VGND VPWR VPWR _07709_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14009_ _06705_ _06706_ _06726_ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__a21oi_1
X_19866_ _01681_ _01689_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__xor2_1
X_18817_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[5\] _11242_ VGND
+ VGND VPWR VPWR _11243_ sky130_fd_sc_hd__xor2_2
XFILLER_0_128_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19797_ top_inst.deskew_buff_inst.col_input\[14\] _11723_ _01622_ _01623_ VGND VGND
+ VPWR VPWR _01624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18748_ _07057_ VGND VGND VPWR VPWR _11177_ sky130_fd_sc_hd__buf_4
XFILLER_0_222_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18679_ net949 _11116_ net167 VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20710_ top_inst.deskew_buff_inst.col_input\[46\] _11723_ _02487_ _02488_ VGND VGND
+ VPWR VPWR _02489_ sky130_fd_sc_hd__a22o_1
XFILLER_0_231_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21690_ _03402_ _03417_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_1322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20641_ _01819_ _02420_ _02421_ _02035_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23360_ net461 _04791_ _04798_ _04795_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20572_ _02316_ _02319_ net175 _02353_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_50_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22311_ _03995_ _03997_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23291_ net743 _04752_ _04759_ _04756_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22242_ _03923_ _03925_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22173_ _03861_ _03862_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21124_ top_inst.grid_inst.data_path_wires\[17\]\[7\] VGND VGND VPWR VPWR _02878_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21055_ _02818_ _02819_ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_219_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20006_ _01815_ _01821_ _01822_ _01820_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__a22o_1
XFILLER_0_185_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21957_ _03655_ _03669_ _03670_ _03654_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__nand4b_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ _02651_ _02665_ _02677_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__and3_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12690_ _05499_ _05500_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_171_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21888_ _03587_ _03605_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__nand2_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23627_ clknet_leaf_100_clk _00160_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20839_ _02594_ _02611_ _07595_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14360_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _07066_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23558_ clknet_leaf_102_clk net915 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13311_ _06083_ _06084_ _06085_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22509_ _04173_ _04161_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__and2b_1
XFILLER_0_135_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput19 input_tdata[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14291_ _06966_ _07000_ VGND VGND VPWR VPWR _07001_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23489_ clknet_leaf_140_clk net615 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[79\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_892 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13242_ _05980_ _06018_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16030_ _08636_ _08637_ VGND VGND VPWR VPWR _08638_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_220_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13173_ _05949_ _05951_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__nor2_1
XFILLER_0_206_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12124_ net793 _05084_ _05085_ _05075_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17981_ net1011 _10364_ _10483_ _10484_ _09886_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19720_ _01546_ _01547_ _01500_ _01523_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__o211ai_2
X_16932_ _09485_ _09486_ _09457_ VGND VGND VPWR VPWR _09488_ sky130_fd_sc_hd__a21o_1
X_12055_ net997 _05045_ _05046_ _05035_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__o211a_1
X_19651_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[11\] _01480_ VGND
+ VGND VPWR VPWR _01481_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_217_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16863_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[8\] _09419_ VGND
+ VGND VPWR VPWR _09420_ sky130_fd_sc_hd__xnor2_1
X_18602_ _11043_ _11061_ VGND VGND VPWR VPWR _11062_ sky130_fd_sc_hd__or2b_1
X_15814_ _08385_ _08386_ _08427_ VGND VGND VPWR VPWR _08428_ sky130_fd_sc_hd__o21a_1
X_19582_ _01410_ _01411_ _01412_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_204_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16794_ _09287_ _09318_ _09350_ _09351_ VGND VGND VPWR VPWR _09353_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18533_ _10961_ _10962_ _10994_ VGND VGND VPWR VPWR _10995_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_232_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15745_ _08357_ _08359_ VGND VGND VPWR VPWR _08360_ sky130_fd_sc_hd__xnor2_2
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12957_ top_inst.grid_inst.data_path_wires\[1\]\[7\] VGND VGND VPWR VPWR _05753_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_834 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11908_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[29\] _04956_
+ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__or2_1
X_18464_ _10925_ _10926_ VGND VGND VPWR VPWR _10927_ sky130_fd_sc_hd__and2b_1
XFILLER_0_201_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15676_ _08283_ _08292_ VGND VGND VPWR VPWR _08293_ sky130_fd_sc_hd__nand2_1
X_12888_ _05664_ _05667_ _05693_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__or3_1
XFILLER_0_158_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17415_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[27\] _09631_ VGND
+ VGND VPWR VPWR _09953_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14627_ _07282_ _07277_ VGND VGND VPWR VPWR _07317_ sky130_fd_sc_hd__or2b_1
XFILLER_0_184_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18395_ _10855_ _10859_ VGND VGND VPWR VPWR _10860_ sky130_fd_sc_hd__xnor2_1
X_11839_ top_inst.axis_out_inst.out_buff_data\[95\] _04917_ VGND VGND VPWR VPWR _04923_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17346_ _09863_ _09883_ VGND VGND VPWR VPWR _09887_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14558_ _07247_ _07248_ _07240_ VGND VGND VPWR VPWR _07250_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13509_ _06240_ _06258_ _05315_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__o21a_1
X_17277_ _09807_ _09821_ VGND VGND VPWR VPWR _09822_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14489_ net171 _07181_ _07182_ VGND VGND VPWR VPWR _07183_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_141_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19016_ _11401_ _11408_ VGND VGND VPWR VPWR _11437_ sky130_fd_sc_hd__or2b_1
XFILLER_0_114_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16228_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[6\] _08811_ VGND
+ VGND VPWR VPWR _08812_ sky130_fd_sc_hd__xor2_2
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16159_ _08743_ _08744_ VGND VGND VPWR VPWR _08745_ sky130_fd_sc_hd__nand2_1
XFILLER_0_228_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_1124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19918_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[20\] _01480_ VGND
+ VGND VPWR VPWR _01739_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_242_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19849_ _01652_ _01673_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__nand2_1
XFILLER_0_236_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22860_ net1043 _04509_ _04512_ _04511_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__o211a_1
XFILLER_0_218_1053 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21811_ _03531_ _03532_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22791_ _04425_ _04421_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24530_ clknet_leaf_129_clk _01063_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_52_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21742_ _03433_ _03436_ VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24461_ clknet_leaf_55_clk _00994_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_21673_ _03070_ _03400_ _03401_ _02909_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23412_ net619 _04596_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20624_ _02001_ _02227_ _02404_ _02186_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__a22o_1
X_24392_ clknet_leaf_39_clk net709 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23343_ net781 _04778_ _04788_ _04782_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20555_ _02297_ _02299_ _02337_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__a21o_1
XFILLER_0_190_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23274_ net377 _04739_ _04749_ _04743_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20486_ _02226_ _02235_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__or2b_1
XFILLER_0_61_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22225_ _03911_ _03913_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_929 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_203_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_242_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22156_ _03846_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21107_ top_inst.grid_inst.data_path_wires\[17\]\[2\] VGND VGND VPWR VPWR _02866_
+ sky130_fd_sc_hd__clkbuf_4
X_22087_ _03709_ _03680_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21038_ _06178_ _02803_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_233_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13860_ _06555_ _06574_ _06572_ VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_198_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12811_ _05614_ _05618_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__and2_1
XFILLER_0_241_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22989_ net965 _04575_ _04585_ _04577_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13791_ _06496_ _06533_ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _08159_ sky130_fd_sc_hd__buf_4
X_12742_ _05525_ _05526_ _05550_ _05551_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__a211oi_4
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12673_ _05468_ _05462_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__or2b_1
X_15461_ _07956_ _08072_ VGND VGND VPWR VPWR _08102_ sky130_fd_sc_hd__and2b_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17200_ _09739_ _09723_ VGND VGND VPWR VPWR _09748_ sky130_fd_sc_hd__or2b_1
X_14412_ _07107_ _07108_ VGND VGND VPWR VPWR _07109_ sky130_fd_sc_hd__xnor2_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18180_ _10648_ _10649_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[3\]
+ VGND VGND VPWR VPWR _10651_ sky130_fd_sc_hd__a21oi_1
X_15392_ _07990_ _08034_ VGND VGND VPWR VPWR _08035_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17131_ _09634_ _09646_ _09645_ VGND VGND VPWR VPWR _09682_ sky130_fd_sc_hd__a21boi_1
X_14343_ _06936_ _07030_ VGND VGND VPWR VPWR _07051_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17062_ _09585_ _09614_ VGND VGND VPWR VPWR _09615_ sky130_fd_sc_hd__xnor2_1
X_14274_ _06945_ _06984_ VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13225_ _05968_ _05963_ _06001_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16013_ _08620_ _08621_ VGND VGND VPWR VPWR _08622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_221_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13156_ top_inst.grid_inst.data_path_wires\[1\]\[4\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[1\]\[5\]
+ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _05009_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__buf_2
XFILLER_0_85_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _05864_ _05867_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__and2_1
X_17964_ _10377_ _10466_ VGND VGND VPWR VPWR _10468_ sky130_fd_sc_hd__or2_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19703_ _01489_ _01491_ _01490_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__a21bo_1
X_16915_ _09360_ _09377_ _09196_ _09201_ VGND VGND VPWR VPWR _09471_ sky130_fd_sc_hd__or4b_4
XFILLER_0_178_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12038_ net262 _05036_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__or2_1
XFILLER_0_236_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17895_ _10357_ _10360_ _10400_ VGND VGND VPWR VPWR _10401_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19634_ _01462_ _01463_ _01422_ _01424_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__o211a_1
X_16846_ _09354_ _09356_ _09352_ VGND VGND VPWR VPWR _09404_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_75_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19565_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[8\] _01395_ _01396_
+ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__a21o_1
X_16777_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[2\] _09206_ _09333_
+ _09334_ VGND VGND VPWR VPWR _09336_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13989_ _06690_ _06695_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__or2b_1
XFILLER_0_177_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1095 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18516_ _10592_ _10612_ _10976_ VGND VGND VPWR VPWR _10978_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_220_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15728_ _08342_ _08343_ VGND VGND VPWR VPWR _08344_ sky130_fd_sc_hd__nor2_1
X_19496_ net197 _01268_ _01328_ _01329_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_87_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_1094 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18447_ _10882_ _10883_ _10910_ VGND VGND VPWR VPWR _10911_ sky130_fd_sc_hd__a21o_1
X_15659_ _08274_ _08275_ VGND VGND VPWR VPWR _08276_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18378_ _10798_ _10800_ _10842_ VGND VGND VPWR VPWR _10843_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17329_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[21\] _09628_ _09629_
+ VGND VGND VPWR VPWR _09871_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20340_ _02092_ _02093_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20271_ _02059_ _02060_ _02041_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22010_ _03709_ _05275_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23961_ clknet_leaf_89_clk _00494_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_192_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22912_ net413 _04535_ _04541_ _04537_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23892_ clknet_leaf_62_clk _00425_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22843_ net674 _04496_ _04502_ _04498_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22774_ net724 _05317_ _04442_ _04443_ _09806_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24513_ clknet_leaf_132_clk _01046_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dfxtp_1
X_21725_ _03449_ _03450_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__nor2_1
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24444_ clknet_leaf_64_clk net980 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[0\].output_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21656_ _03356_ _03373_ _03383_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__and3_1
XFILLER_0_192_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20607_ _02215_ _02220_ _02386_ _02384_ _02387_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__o41a_1
XFILLER_0_227_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24375_ clknet_leaf_39_clk net395 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].output_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21587_ _03246_ _03316_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23326_ _04686_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__buf_4
XFILLER_0_104_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20538_ _02319_ net176 VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_1280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23257_ _04686_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20469_ _02251_ _02252_ _02236_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__a21o_1
X_13010_ _05741_ _05759_ _05757_ _05744_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22208_ _03889_ _03896_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__xnor2_2
XTAP_6600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23188_ _04686_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__buf_2
XTAP_6611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22139_ _03824_ _03829_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__xnor2_1
XTAP_6644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14961_ _07624_ _07611_ _07625_ _07618_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__o211a_1
XTAP_6699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16700_ _09243_ _09261_ VGND VGND VPWR VPWR _09262_ sky130_fd_sc_hd__or2_2
X_13912_ _06640_ _06641_ VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__or2_1
XTAP_5987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17680_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[6\] _10190_ _08307_
+ VGND VGND VPWR VPWR _10191_ sky130_fd_sc_hd__mux2_1
XTAP_5998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14892_ net1088 _07048_ _07574_ _07575_ _06180_ VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__o221a_1
XFILLER_0_230_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16631_ top_inst.skew_buff_inst.row\[2\].output_reg\[3\] top_inst.axis_in_inst.inbuf_bus\[19\]
+ _07059_ VGND VGND VPWR VPWR _09201_ sky130_fd_sc_hd__mux2_4
X_13843_ _06364_ _06584_ VGND VGND VPWR VPWR _06585_ sky130_fd_sc_hd__and2_1
XFILLER_0_242_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19350_ _11684_ _11679_ _11687_ _11692_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__nand4_1
XFILLER_0_187_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16562_ _09103_ _09104_ VGND VGND VPWR VPWR _09138_ sky130_fd_sc_hd__or2b_1
XFILLER_0_69_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13774_ _06515_ _06517_ VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18301_ top_inst.grid_inst.data_path_wires\[12\]\[1\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _10768_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15513_ top_inst.grid_inst.data_path_wires\[7\]\[5\] VGND VGND VPWR VPWR _08147_
+ sky130_fd_sc_hd__buf_4
XFILLER_0_231_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12725_ _05293_ _05297_ _05301_ _05288_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__a22oi_2
X_19281_ _11683_ VGND VGND VPWR VPWR _11684_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_155_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_242_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16493_ _09069_ _09070_ VGND VGND VPWR VPWR _09071_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18232_ _10646_ _10667_ VGND VGND VPWR VPWR _10701_ sky130_fd_sc_hd__nor2_1
X_15444_ _08084_ _08085_ VGND VGND VPWR VPWR _08086_ sky130_fd_sc_hd__nand2_1
XFILLER_0_242_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12656_ _05466_ _05467_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18163_ _10628_ _10634_ VGND VGND VPWR VPWR _10635_ sky130_fd_sc_hd__or2_1
X_12587_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[5\] _05354_ _05398_
+ _05400_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15375_ _08016_ _08018_ VGND VGND VPWR VPWR _08019_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_974 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17114_ _09654_ _09655_ _09653_ VGND VGND VPWR VPWR _09665_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14326_ _06980_ _07034_ VGND VGND VPWR VPWR _07035_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18094_ _10581_ _08674_ VGND VGND VPWR VPWR _10582_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold408 top_inst.axis_in_inst.inbuf_bus\[20\] VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17045_ _09361_ _09377_ _09210_ _09214_ VGND VGND VPWR VPWR _09598_ sky130_fd_sc_hd__or4b_4
Xhold419 _00235_ VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__dlygate4sd3_1
X_14257_ _06964_ _06965_ VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13208_ _05982_ _05985_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_1239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14188_ _06860_ _06900_ VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__xnor2_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13139_ _05916_ _05918_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18996_ _11362_ _11364_ VGND VGND VPWR VPWR _11418_ sky130_fd_sc_hd__nor2_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17947_ _10411_ _10417_ _10415_ VGND VGND VPWR VPWR _10451_ sky130_fd_sc_hd__a21o_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17878_ _10381_ _10383_ VGND VGND VPWR VPWR _10384_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_233_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16829_ _09384_ _09385_ _09370_ VGND VGND VPWR VPWR _09387_ sky130_fd_sc_hd__a21o_1
X_19617_ _01445_ _01446_ _01447_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__nand3_1
XFILLER_0_221_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19548_ _01349_ _01380_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__xor2_2
XFILLER_0_221_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19479_ _11701_ net248 VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21510_ _03201_ _03204_ _03242_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_152_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22490_ _04132_ _04144_ _04171_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21441_ _03172_ _03175_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24160_ clknet_leaf_9_clk _00693_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21372_ _03105_ _03108_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_160_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23111_ top_inst.axis_out_inst.out_buff_enabled _04857_ VGND VGND VPWR VPWR _04654_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20323_ top_inst.grid_inst.data_path_wires\[16\]\[3\] _01992_ _02013_ _02051_ VGND
+ VGND VPWR VPWR _02111_ sky130_fd_sc_hd__nand4_1
X_24091_ clknet_leaf_97_clk _00624_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold920 top_inst.deskew_buff_inst.col_input\[63\] VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold931 top_inst.axis_in_inst.inbuf_bus\[31\] VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__dlygate4sd3_1
X_23042_ net969 _04616_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20254_ _10083_ _02043_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_229_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20185_ top_inst.grid_inst.data_path_wires\[16\]\[2\] VGND VGND VPWR VPWR _01992_
+ sky130_fd_sc_hd__buf_2
XFILLER_0_110_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23944_ clknet_leaf_91_clk _00477_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23875_ clknet_leaf_51_clk _00408_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_233_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22826_ _04490_ _04491_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_233_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22757_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[27\] _04163_ VGND
+ VGND VPWR VPWR _04427_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12510_ _05327_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__buf_8
XFILLER_0_164_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13490_ net1031 _05788_ _06241_ _06207_ VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21708_ _03433_ _03434_ VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__and2_1
X_22688_ _04301_ _04322_ _04360_ _04357_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__and4_1
XFILLER_0_87_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12441_ _05267_ _04863_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24427_ clknet_leaf_54_clk net773 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].output_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21639_ net544 _05316_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__or2_1
XFILLER_0_191_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15160_ _07768_ _07769_ VGND VGND VPWR VPWR _07809_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12372_ net398 _05222_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24358_ clknet_4_5__leaf_clk _00891_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[117\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_244_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14111_ _06785_ _06825_ VGND VGND VPWR VPWR _06826_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15091_ _07710_ _07728_ VGND VGND VPWR VPWR _07741_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23309_ net146 _04766_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_240_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24289_ clknet_leaf_12_clk _00822_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14042_ _06735_ _06736_ _06757_ VGND VGND VPWR VPWR _06759_ sky130_fd_sc_hd__and3_1
XFILLER_0_240_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18850_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[13\]\[3\]
+ top_inst.grid_inst.data_path_wires\[13\]\[2\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[4\]
+ VGND VGND VPWR VPWR _11275_ sky130_fd_sc_hd__a22oi_1
XTAP_6430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17801_ _10307_ _10308_ VGND VGND VPWR VPWR _10309_ sky130_fd_sc_hd__nor2_1
XFILLER_0_234_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18781_ _10641_ _11208_ VGND VGND VPWR VPWR _11209_ sky130_fd_sc_hd__and2_1
XTAP_6485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15993_ _08600_ _08601_ VGND VGND VPWR VPWR _08602_ sky130_fd_sc_hd__or2b_1
XTAP_5751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17732_ _10035_ _10032_ _10052_ _10050_ VGND VGND VPWR VPWR _10241_ sky130_fd_sc_hd__nand4_2
XTAP_5773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14944_ top_inst.grid_inst.data_path_wires\[6\]\[3\] VGND VGND VPWR VPWR _07613_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17663_ _10032_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[2\] _10171_
+ _10172_ VGND VGND VPWR VPWR _10174_ sky130_fd_sc_hd__o2bb2a_1
X_14875_ _07521_ _07525_ _07523_ VGND VGND VPWR VPWR _07559_ sky130_fd_sc_hd__a21o_1
XFILLER_0_202_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19402_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[4\] net192 net247
+ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _01238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16614_ _09186_ VGND VGND VPWR VPWR _09187_ sky130_fd_sc_hd__buf_2
XFILLER_0_159_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13826_ _06532_ _06531_ VGND VGND VPWR VPWR _06568_ sky130_fd_sc_hd__or2b_1
X_17594_ top_inst.grid_inst.data_path_wires\[11\]\[3\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[11\]\[4\]
+ VGND VGND VPWR VPWR _10107_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_724 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19333_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[2\] _11725_ _11726_
+ VGND VGND VPWR VPWR _11727_ sky130_fd_sc_hd__nand3_1
XFILLER_0_187_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16545_ _09118_ _09119_ _09040_ _09120_ VGND VGND VPWR VPWR _09121_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13757_ _06456_ _06455_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_136_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_136_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_134_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12708_ _05516_ _05517_ _05484_ _05485_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__o211a_1
X_19264_ net959 _11662_ _11675_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16476_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[11\] _08975_ _08896_
+ VGND VGND VPWR VPWR _09054_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13688_ _06382_ _06380_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_667 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18215_ _10577_ _10610_ VGND VGND VPWR VPWR _10684_ sky130_fd_sc_hd__nand2_1
X_15427_ _07624_ _07640_ _07637_ VGND VGND VPWR VPWR _08069_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_1396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12639_ _05448_ _05450_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__nand2_1
X_19195_ _11575_ _11550_ VGND VGND VPWR VPWR _11612_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18146_ _10447_ VGND VGND VPWR VPWR _10620_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15358_ _07989_ _07965_ _08000_ VGND VGND VPWR VPWR _08002_ sky130_fd_sc_hd__nand3_1
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold205 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[2\] VGND VGND
+ VPWR VPWR net387 sky130_fd_sc_hd__dlygate4sd3_1
X_14309_ _07015_ _07017_ VGND VGND VPWR VPWR _07019_ sky130_fd_sc_hd__and2_1
XFILLER_0_170_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18077_ net946 _10563_ _10576_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__o21a_1
XFILLER_0_223_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15289_ _07933_ _07934_ VGND VGND VPWR VPWR _07935_ sky130_fd_sc_hd__xnor2_2
Xhold216 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[4\] VGND
+ VGND VPWR VPWR net398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold227 _00201_ VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 top_inst.deskew_buff_inst.col_input\[11\] VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ _09529_ VGND VGND VPWR VPWR _09581_ sky130_fd_sc_hd__inv_2
Xhold249 _00065_ VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18979_ _11399_ _11400_ VGND VGND VPWR VPWR _11401_ sky130_fd_sc_hd__xor2_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21990_ _03695_ _03691_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__or2_1
X_20941_ _02635_ _02709_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__and2b_1
XFILLER_0_234_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23660_ clknet_leaf_135_clk _00193_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_20872_ _02643_ _02622_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22611_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[19\] _04215_ _04216_
+ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23591_ clknet_leaf_101_clk _00124_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_127_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_127_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22542_ _04220_ _04221_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__and2b_1
XFILLER_0_130_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_976 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22473_ _04152_ _04155_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21424_ net924 _02491_ _03158_ _03159_ _02962_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__o221a_1
X_24212_ clknet_leaf_118_clk _00745_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24143_ clknet_leaf_18_clk _00676_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_114_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21355_ _03090_ _03091_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_142_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_241_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_999 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20306_ _02050_ _02067_ _02066_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__o21ba_1
X_24074_ clknet_leaf_112_clk _00607_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21286_ _03022_ _03023_ _02993_ _02994_ VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__o211ai_1
Xhold750 top_inst.deskew_buff_inst.col_input\[1\] VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[15\] VGND
+ VGND VPWR VPWR net943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23025_ net23 _04601_ _04607_ _04606_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__o211a_1
Xhold772 top_inst.deskew_buff_inst.col_input\[95\] VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__buf_1
Xhold783 top_inst.axis_in_inst.inbuf_bus\[12\] VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__dlygate4sd3_1
X_20237_ _02007_ _02028_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold794 top_inst.deskew_buff_inst.col_input\[25\] VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__buf_1
XFILLER_0_228_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20168_ _01563_ _01977_ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__xnor2_1
XTAP_5036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_239_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20099_ _01824_ _01909_ _01911_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__a21o_1
X_12990_ net1044 _05314_ _05776_ _05767_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__o211a_1
XTAP_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23927_ clknet_leaf_76_clk _00460_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _04874_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_1042 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _07318_ _07349_ VGND VGND VPWR VPWR _07350_ sky130_fd_sc_hd__xnor2_4
XTAP_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23858_ clknet_leaf_77_clk _00391_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _04874_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__buf_2
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _06320_ _06322_ _06358_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__or3_1
XFILLER_0_184_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22809_ net666 _09804_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14591_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[8\] _07281_ VGND
+ VGND VPWR VPWR _07282_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_118_clk clknet_4_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23789_ clknet_leaf_70_clk _00322_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_156_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16330_ _08855_ _08856_ _08911_ VGND VGND VPWR VPWR _08912_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13542_ _06271_ _06276_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16261_ _08838_ _08843_ VGND VGND VPWR VPWR _08844_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13473_ _06181_ _06205_ _06225_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18000_ _10377_ _10502_ VGND VGND VPWR VPWR _10503_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_164_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15212_ _07803_ _07804_ _07859_ VGND VGND VPWR VPWR _07860_ sky130_fd_sc_hd__a21oi_1
X_12424_ _05177_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__clkbuf_8
X_16192_ _08772_ _08776_ VGND VGND VPWR VPWR _08777_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15143_ _07786_ _07791_ VGND VGND VPWR VPWR _07792_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12355_ _05177_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_239_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19951_ _01769_ _01770_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__xor2_2
X_15074_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[5\] _07724_ VGND
+ VGND VPWR VPWR _07725_ sky130_fd_sc_hd__xor2_2
XFILLER_0_121_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12286_ _05177_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14025_ _06740_ _06741_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__nand2_1
X_18902_ _11324_ _11325_ VGND VGND VPWR VPWR _11326_ sky130_fd_sc_hd__xnor2_1
X_19882_ _01663_ _01664_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18833_ _11230_ _11246_ VGND VGND VPWR VPWR _11258_ sky130_fd_sc_hd__nand2_1
XTAP_6260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18764_ _11154_ _11132_ _11130_ _11156_ VGND VGND VPWR VPWR _11192_ sky130_fd_sc_hd__a22o_1
XTAP_5570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15976_ _08582_ _08584_ VGND VGND VPWR VPWR _08586_ sky130_fd_sc_hd__or2_1
XFILLER_0_234_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17715_ _10187_ _10189_ _10186_ VGND VGND VPWR VPWR _10225_ sky130_fd_sc_hd__o21bai_2
X_14927_ _07593_ _07602_ _07594_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__o21a_1
X_18695_ _11138_ _11133_ VGND VGND VPWR VPWR _11139_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17646_ _10134_ _10140_ VGND VGND VPWR VPWR _10157_ sky130_fd_sc_hd__or2b_1
X_14858_ _07487_ _07491_ _07489_ VGND VGND VPWR VPWR _07543_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13809_ _06522_ _06519_ _06550_ _06404_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__a31oi_1
X_17577_ _10027_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[0\]
+ _10029_ VGND VGND VPWR VPWR _10091_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_109_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_16
X_14789_ _07473_ _07474_ _07448_ VGND VGND VPWR VPWR _07476_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_202_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19316_ _11679_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[0\] _11677_
+ VGND VGND VPWR VPWR _11712_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16528_ _09103_ _09104_ VGND VGND VPWR VPWR _09105_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19247_ _11177_ _11660_ _11661_ _11641_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16459_ _08999_ _09037_ _05335_ VGND VGND VPWR VPWR _09038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19178_ _11589_ _11593_ VGND VGND VPWR VPWR _11595_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18129_ _05755_ VGND VGND VPWR VPWR _10607_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_223_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21140_ _02889_ _02021_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21071_ _02818_ _02819_ _02816_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__o21a_1
XFILLER_0_158_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20022_ net786 _01386_ VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__or2_1
XFILLER_0_226_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1015 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21973_ top_inst.grid_inst.data_path_wires\[18\]\[2\] VGND VGND VPWR VPWR _03684_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_193_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer20 _09214_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer31 net211 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__buf_1
XFILLER_0_154_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer42 _09196_ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__buf_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23712_ clknet_leaf_123_clk _00245_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer53 _11699_ VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_1
X_20924_ _02518_ _02693_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer64 _11686_ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer75 _07081_ VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23643_ clknet_leaf_126_clk net374 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_20855_ _02626_ _02627_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23574_ clknet_leaf_108_clk net498 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_20786_ _02527_ _02547_ _02561_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22525_ _04189_ _04190_ _04204_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__or3_1
XFILLER_0_106_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22456_ _03693_ _04138_ _04102_ _04104_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21407_ _02868_ _02893_ _03092_ _03142_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__a31o_1
X_22387_ _03711_ _03690_ _04027_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12140_ net930 _05084_ _05094_ _05088_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__o211a_1
XFILLER_0_241_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24126_ clknet_leaf_118_clk _00659_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_21338_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[7\] _03038_ _03039_
+ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_103_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12071_ net556 _05045_ _05055_ _05049_ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__o211a_1
X_24057_ clknet_leaf_46_clk _00590_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_21269_ _02862_ _02895_ _02893_ _02864_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__a22oi_1
Xhold580 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[0\]\[1\] VGND VGND
+ VPWR VPWR net762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold591 _00960_ VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23008_ _04863_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_216_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ _08441_ _08442_ VGND VGND VPWR VPWR _08443_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _08318_ _08320_ _08375_ VGND VGND VPWR VPWR _08376_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_204_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12973_ _05744_ _05756_ _05764_ _05743_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__o211a_1
XFILLER_0_232_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17500_ _04858_ VGND VGND VPWR VPWR _10030_ sky130_fd_sc_hd__buf_2
XTAP_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14712_ _07359_ _07400_ VGND VGND VPWR VPWR _07401_ sky130_fd_sc_hd__xnor2_1
XTAP_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ _10901_ _10900_ VGND VGND VPWR VPWR _10943_ sky130_fd_sc_hd__or2b_1
X_11924_ net478 _04964_ _04971_ _04968_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__o211a_1
XTAP_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _08197_ _08308_ VGND VGND VPWR VPWR _08309_ sky130_fd_sc_hd__and2_1
XFILLER_0_231_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17431_ _09932_ _09946_ _09968_ VGND VGND VPWR VPWR _09969_ sky130_fd_sc_hd__a21oi_1
XTAP_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _07072_ VGND VGND VPWR VPWR _07333_ sky130_fd_sc_hd__inv_2
XFILLER_0_197_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11855_ net921 _04925_ _04932_ _04929_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__o211a_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17362_ _09872_ _09878_ _09900_ _09855_ VGND VGND VPWR VPWR _09903_ sky130_fd_sc_hd__a22o_1
XFILLER_0_184_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14574_ _07263_ _07264_ _07217_ VGND VGND VPWR VPWR _07266_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11786_ net757 _04890_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__or2_1
X_19101_ _11147_ _11161_ VGND VGND VPWR VPWR _11520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16313_ top_inst.grid_inst.data_path_wires\[8\]\[7\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _08895_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13525_ _06273_ _06274_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__nor2_1
X_17293_ _09624_ _09835_ VGND VGND VPWR VPWR _09837_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19032_ _11435_ _11452_ VGND VGND VPWR VPWR _11453_ sky130_fd_sc_hd__xnor2_1
X_16244_ _08826_ _08827_ VGND VGND VPWR VPWR _08828_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13456_ _06193_ _06204_ _06213_ _06207_ VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12407_ _05127_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__buf_2
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16175_ _08758_ _08759_ _07057_ VGND VGND VPWR VPWR _08761_ sky130_fd_sc_hd__a21o_1
X_13387_ _06113_ _06132_ _06130_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__a21oi_1
Xoutput107 net107 VGND VGND VPWR VPWR output_tdata[47] sky130_fd_sc_hd__buf_2
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput118 net118 VGND VGND VPWR VPWR output_tdata[57] sky130_fd_sc_hd__clkbuf_4
X_15126_ _07681_ _07703_ _07732_ _07736_ VGND VGND VPWR VPWR _07776_ sky130_fd_sc_hd__o31a_1
Xoutput129 net129 VGND VGND VPWR VPWR output_tdata[67] sky130_fd_sc_hd__buf_2
XFILLER_0_50_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12338_ _05127_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__buf_2
XFILLER_0_239_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19934_ _01749_ _01754_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__nand2_1
X_15057_ net1071 _07048_ _07705_ _07706_ _07708_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__o221a_1
XFILLER_0_120_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12269_ net934 _05164_ _05167_ _05168_ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14008_ _06723_ _06725_ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_177_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19865_ _01665_ _01688_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_235_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18816_ _11240_ _11241_ VGND VGND VPWR VPWR _11242_ sky130_fd_sc_hd__nand2_1
XTAP_6090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19796_ _01621_ _01594_ _01595_ _05311_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__o31a_1
XFILLER_0_235_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15959_ _08557_ _08525_ _08567_ VGND VGND VPWR VPWR _08569_ sky130_fd_sc_hd__nand3_1
X_18747_ net977 _10616_ _11176_ _11160_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18678_ net1009 _11116_ net167 VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__o21a_1
XFILLER_0_210_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17629_ _10134_ _10140_ VGND VGND VPWR VPWR _10141_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20640_ net816 _01386_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__or2_1
XFILLER_0_191_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20571_ _02315_ _02322_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22310_ _03951_ _03959_ _03996_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23290_ net137 _04753_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22241_ _03070_ _03927_ _03928_ _03929_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22172_ _03707_ _03688_ _03705_ _03686_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__nand4_1
XFILLER_0_160_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21123_ _10583_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_2_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21054_ _02674_ _02788_ _02791_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20005_ _01753_ _01793_ _01794_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__a21o_1
XFILLER_0_201_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_1002 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21956_ _03665_ _03652_ _03668_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__nand3_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _02651_ _02665_ _02677_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__a21oi_2
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21887_ _03587_ _03605_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__or2_1
XFILLER_0_171_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23626_ clknet_leaf_100_clk net386 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_20838_ _02594_ _02611_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23557_ clknet_leaf_102_clk _00090_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20769_ _01819_ _02544_ _02545_ _02035_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__o211a_1
X_13310_ _05753_ _05768_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__nand2_1
X_22508_ _04170_ _04172_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__nor2_1
X_14290_ _06998_ _06999_ VGND VGND VPWR VPWR _07000_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23488_ clknet_leaf_140_clk net571 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[78\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13241_ _05751_ _06016_ _06017_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__a21oi_1
X_22439_ net627 _09804_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13172_ _05947_ _05948_ _05950_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_27_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24109_ clknet_leaf_16_clk _00642_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12123_ net791 _05076_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17980_ _10449_ _10443_ _10482_ _07439_ VGND VGND VPWR VPWR _10484_ sky130_fd_sc_hd__a31o_1
XFILLER_0_237_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16931_ _09457_ _09485_ _09486_ VGND VGND VPWR VPWR _09487_ sky130_fd_sc_hd__nand3_1
X_12054_ net256 _05036_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__or2_1
XFILLER_0_217_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16862_ _09418_ _09417_ VGND VGND VPWR VPWR _09419_ sky130_fd_sc_hd__nor2_8
X_19650_ _01354_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__buf_4
XFILLER_0_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18601_ _11051_ _11060_ VGND VGND VPWR VPWR _11061_ sky130_fd_sc_hd__xnor2_1
X_15813_ _08382_ _08384_ VGND VGND VPWR VPWR _08427_ sky130_fd_sc_hd__or2_1
XFILLER_0_232_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19581_ _01410_ _01411_ _01412_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__nand3_1
XFILLER_0_244_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16793_ _09287_ _09318_ _09350_ _09351_ VGND VGND VPWR VPWR _09352_ sky130_fd_sc_hd__or4_1
XFILLER_0_137_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18532_ _10964_ _10993_ VGND VGND VPWR VPWR _10994_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15744_ _08311_ _08312_ _08358_ VGND VGND VPWR VPWR _08359_ sky130_fd_sc_hd__o21ba_1
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12956_ _05751_ _05735_ _05752_ _05743_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11907_ net668 _04951_ _04961_ _04955_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _10595_ _10602_ _10893_ _10892_ _10592_ VGND VGND VPWR VPWR _10926_ sky130_fd_sc_hd__a32o_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ _08284_ _08291_ VGND VGND VPWR VPWR _08292_ sky130_fd_sc_hd__xnor2_1
X_12887_ _05691_ _05692_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__and2_1
XFILLER_0_158_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_975 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17414_ _09915_ _09935_ _09913_ VGND VGND VPWR VPWR _09952_ sky130_fd_sc_hd__o21a_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _07308_ _07309_ _07315_ VGND VGND VPWR VPWR _07316_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18394_ _10856_ _10858_ VGND VGND VPWR VPWR _10859_ sky130_fd_sc_hd__nor2_1
X_11838_ net689 _04912_ _04922_ _04916_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17345_ net1047 _09266_ _09884_ _09885_ _09886_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14557_ _07240_ _07247_ _07248_ VGND VGND VPWR VPWR _07249_ sky130_fd_sc_hd__nand3_1
XFILLER_0_126_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11769_ net622 _04877_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_184_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13508_ _06240_ _06258_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__nand2_1
X_17276_ _09819_ _09820_ VGND VGND VPWR VPWR _09821_ sky130_fd_sc_hd__and2_1
X_14488_ _07140_ _07143_ VGND VGND VPWR VPWR _07182_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19015_ _11407_ _11406_ VGND VGND VPWR VPWR _11436_ sky130_fd_sc_hd__or2b_1
X_16227_ _08809_ _08810_ VGND VGND VPWR VPWR _08811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13439_ _06181_ _05756_ _06201_ _06183_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16158_ _08671_ _08669_ _08686_ _08682_ VGND VGND VPWR VPWR _08744_ sky130_fd_sc_hd__nand4_1
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15109_ _07756_ _07757_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[6\]
+ VGND VGND VPWR VPWR _07759_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16089_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _08686_ sky130_fd_sc_hd__buf_2
XFILLER_0_227_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1081 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19917_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[19\] _01395_ _01396_
+ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__a21o_2
XFILLER_0_227_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1013 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19848_ _01671_ _01672_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__and2_1
XFILLER_0_235_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19779_ _11703_ _11709_ _01534_ _01605_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__a211o_2
X_21810_ _03278_ _03530_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22790_ _04407_ _04458_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21741_ _03438_ _03463_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__nand2_1
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24460_ clknet_leaf_55_clk _00993_ VGND VGND VPWR VPWR top_inst.axis_in_inst.inbuf_bus\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21672_ net411 _02638_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__or2_1
XFILLER_0_231_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23411_ net467 _04856_ _04870_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__o21a_1
XFILLER_0_164_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1062 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20623_ _02001_ _02020_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__nand2_1
X_24391_ clknet_leaf_38_clk net295 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_31_clk clknet_4_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23342_ net162 _04779_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20554_ _02323_ _02336_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23273_ net129 _04740_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__or2_1
X_20485_ _02222_ _02259_ VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22224_ _03865_ _03871_ _03912_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__o21a_1
XFILLER_0_203_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22155_ _03311_ _03845_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21106_ _01990_ _11142_ _02865_ _02707_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22086_ _03764_ _03769_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__and2b_1
X_21037_ _02763_ _02783_ _02801_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12810_ _05616_ _05617_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__nor2_1
XFILLER_0_198_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13790_ _06531_ _06532_ VGND VGND VPWR VPWR _06533_ sky130_fd_sc_hd__xnor2_1
X_22988_ net718 _04583_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__or2_1
XFILLER_0_241_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_214_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12741_ _05545_ _05549_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21939_ _03453_ _03617_ _03633_ _03635_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__o31a_1
XFILLER_0_70_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15460_ _08075_ _08082_ _08074_ VGND VGND VPWR VPWR _08101_ sky130_fd_sc_hd__a21oi_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ net1013 _05403_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14411_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[1\] _07096_ _07097_
+ VGND VGND VPWR VPWR _07108_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23609_ clknet_leaf_104_clk net547 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_15391_ _08032_ _08033_ VGND VGND VPWR VPWR _08034_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24589_ clknet_leaf_32_clk _01122_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_22_clk clknet_4_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_231_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17130_ _09670_ _09680_ VGND VGND VPWR VPWR _09681_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_167_1237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14342_ _06979_ _07049_ VGND VGND VPWR VPWR _07050_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_163_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17061_ _09587_ _09613_ VGND VGND VPWR VPWR _09614_ sky130_fd_sc_hd__xor2_1
X_14273_ _06982_ _06983_ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16012_ _08543_ _08545_ _08587_ _08588_ _08590_ VGND VGND VPWR VPWR _08621_ sky130_fd_sc_hd__a32o_2
X_13224_ _05968_ _05963_ _06001_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__a21o_1
XFILLER_0_243_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13155_ _05931_ _05933_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ net501 _05071_ _05074_ _05075_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13086_ _05865_ _05866_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__nor2_1
X_17963_ _10377_ _10466_ VGND VGND VPWR VPWR _10467_ sky130_fd_sc_hd__nand2_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_89_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_16
X_19702_ _01526_ _01530_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16914_ _09211_ _09206_ VGND VGND VPWR VPWR _09470_ sky130_fd_sc_hd__and2_1
X_12037_ _05009_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_109_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17894_ _10354_ _10399_ VGND VGND VPWR VPWR _10400_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19633_ _01422_ _01424_ net238 _01463_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16845_ _09401_ _09402_ VGND VGND VPWR VPWR _09403_ sky130_fd_sc_hd__and2b_1
XFILLER_0_233_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16776_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[2\] _09206_ _09333_
+ _09334_ VGND VGND VPWR VPWR _09335_ sky130_fd_sc_hd__nand4_2
X_19564_ _01353_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__clkbuf_4
X_13988_ _06675_ _06697_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__or2_1
XFILLER_0_220_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15727_ _08303_ _08305_ _08302_ VGND VGND VPWR VPWR _08343_ sky130_fd_sc_hd__o21bai_2
X_18515_ _10591_ _10612_ _10976_ VGND VGND VPWR VPWR _10977_ sky130_fd_sc_hd__and3_1
X_12939_ _05738_ _05735_ _05740_ _05308_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19495_ _01325_ _01326_ _01327_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_238_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15658_ _08137_ top_inst.grid_inst.data_path_wires\[7\]\[0\] _08169_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[5\]
+ VGND VGND VPWR VPWR _08275_ sky130_fd_sc_hd__nand4_2
X_18446_ _10884_ _10909_ VGND VGND VPWR VPWR _10910_ sky130_fd_sc_hd__xor2_1
XFILLER_0_186_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_1383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14609_ _07247_ _07249_ VGND VGND VPWR VPWR _07300_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18377_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[9\] _10793_ VGND
+ VGND VPWR VPWR _10842_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15589_ _08207_ _08208_ VGND VGND VPWR VPWR _08209_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk clknet_4_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17328_ _09839_ _09869_ VGND VGND VPWR VPWR _09870_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17259_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[19\] _09804_ VGND
+ VGND VPWR VPWR _09805_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20270_ _01995_ _02007_ _02056_ _02058_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1067 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23960_ clknet_leaf_89_clk _00493_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_22911_ top_inst.skew_buff_inst.row\[2\].output_reg\[3\] _04530_ VGND VGND VPWR VPWR
+ _04541_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23891_ clknet_leaf_51_clk _00424_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22842_ top_inst.skew_buff_inst.row\[3\].output_reg\[5\] _03691_ VGND VGND VPWR VPWR
+ _04502_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_1196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22773_ _04409_ _04421_ _04441_ _06734_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_1135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24512_ clknet_leaf_135_clk _01045_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_94_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21724_ _03278_ _03448_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24443_ clknet_leaf_63_clk net952 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[0\].output_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21655_ _03356_ _03373_ _03383_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20606_ _02352_ _02350_ _02380_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__o21ai_1
X_24374_ clknet_leaf_40_clk net675 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].output_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21586_ _03246_ _03316_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__nor2_1
XFILLER_0_244_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23325_ _04684_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__buf_4
X_20537_ _01995_ _02229_ _02317_ _02318_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__nor4_1
XFILLER_0_62_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_240_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23256_ _04684_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__buf_4
X_20468_ _02236_ _02251_ _02252_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__nand3_1
XFILLER_0_132_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22207_ _03890_ _03895_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__xor2_2
XFILLER_0_28_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23187_ _04684_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__clkbuf_4
X_20399_ _02137_ _02184_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__xor2_1
XTAP_6601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22138_ _03827_ _03828_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__nor2_1
XTAP_5900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14960_ _05736_ _07090_ VGND VGND VPWR VPWR _07625_ sky130_fd_sc_hd__or2_1
XTAP_6689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22069_ _03740_ _03761_ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__xnor2_2
XTAP_5955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13911_ _05772_ VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__buf_2
XTAP_5977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14891_ _07557_ _07573_ _07057_ VGND VGND VPWR VPWR _07575_ sky130_fd_sc_hd__a21o_1
XTAP_5999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16630_ _09185_ _09197_ _09200_ _09184_ VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13842_ _06581_ _06583_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[13\]
+ _05327_ VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_226_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16561_ _09135_ _09136_ VGND VGND VPWR VPWR _09137_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_230_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13773_ _06430_ _06473_ _06516_ VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__a21oi_1
X_18300_ top_inst.grid_inst.data_path_wires\[12\]\[2\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[5\]
+ VGND VGND VPWR VPWR _10767_ sky130_fd_sc_hd__nand2_1
X_15512_ _07615_ _06634_ _08146_ _08142_ VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12724_ _05532_ _05533_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__xnor2_1
X_19280_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _11683_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16492_ _09066_ _09068_ VGND VGND VPWR VPWR _09070_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_242_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18231_ _10683_ _10699_ VGND VGND VPWR VPWR _10700_ sky130_fd_sc_hd__xor2_2
XFILLER_0_210_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15443_ _08067_ _08049_ _08083_ VGND VGND VPWR VPWR _08085_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12655_ _05463_ _05465_ _05304_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18162_ _10632_ _10633_ VGND VGND VPWR VPWR _10634_ sky130_fd_sc_hd__xor2_1
XFILLER_0_154_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15374_ _07976_ _07977_ _08017_ VGND VGND VPWR VPWR _08018_ sky130_fd_sc_hd__a21bo_1
X_12586_ _05372_ _05397_ _05399_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17113_ _09583_ _09662_ _09663_ VGND VGND VPWR VPWR _09664_ sky130_fd_sc_hd__o21a_1
X_14325_ _07032_ _07033_ VGND VGND VPWR VPWR _07034_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18093_ top_inst.grid_inst.data_path_wires\[12\]\[2\] VGND VGND VPWR VPWR _10581_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold409 _00946_ VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__dlygate4sd3_1
X_17044_ _09596_ VGND VGND VPWR VPWR _09597_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14256_ _06964_ _06965_ _06966_ VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13207_ _05931_ _05983_ _05984_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_238_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14187_ _06632_ _06898_ _06899_ VGND VGND VPWR VPWR _06900_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _05852_ _05917_ _05874_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__a21oi_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _11386_ _11416_ VGND VGND VPWR VPWR _11417_ sky130_fd_sc_hd__xor2_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13069_ _05830_ _05835_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__nand2_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17946_ _10405_ _10406_ _10438_ VGND VGND VPWR VPWR _10450_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_2_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_174_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17877_ _10038_ _10054_ _10379_ _10382_ VGND VGND VPWR VPWR _10383_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_75_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19616_ _01298_ _11691_ _11695_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_117_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16828_ _09370_ _09384_ _09385_ VGND VGND VPWR VPWR _09386_ sky130_fd_sc_hd__nand3_2
XFILLER_0_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19547_ _01378_ _01379_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__nor2_2
XFILLER_0_215_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16759_ _09259_ _09289_ _09287_ VGND VGND VPWR VPWR _09319_ sky130_fd_sc_hd__o21a_1
XFILLER_0_221_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19478_ _01308_ _01311_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18429_ _10591_ _10608_ _10604_ top_inst.grid_inst.data_path_wires\[12\]\[7\] VGND
+ VGND VPWR VPWR _10893_ sky130_fd_sc_hd__a22o_1
XFILLER_0_185_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21440_ _03173_ _03174_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21371_ _03106_ _03107_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__and2_1
XFILLER_0_185_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23110_ net620 _10541_ _04653_ _04643_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__o211a_1
X_20322_ top_inst.grid_inst.data_path_wires\[16\]\[2\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[3\]
+ _02051_ top_inst.grid_inst.data_path_wires\[16\]\[3\] VGND VGND VPWR VPWR _02110_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24090_ clknet_leaf_97_clk _00623_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold910 top_inst.deskew_buff_inst.col_input\[11\] VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold921 top_inst.deskew_buff_inst.col_input\[98\] VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_222_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold932 top_inst.axis_in_inst.inbuf_bus\[27\] VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23041_ _04602_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__buf_2
XFILLER_0_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20253_ _10083_ _02043_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20184_ _01990_ _10033_ _01991_ _01840_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23943_ clknet_leaf_85_clk _00476_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23874_ clknet_leaf_50_clk _00407_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22825_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[31\] _04483_ VGND
+ VGND VPWR VPWR _04491_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_233_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22756_ _04390_ _04410_ _04388_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsplit47 _07593_ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_137_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21707_ _03431_ _03432_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__or2_1
X_22687_ _04339_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24426_ clknet_leaf_58_clk net603 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].output_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12440_ net211 VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21638_ _03347_ _03343_ _03366_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__and3_1
XFILLER_0_168_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24357_ clknet_leaf_22_clk _00890_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[116\]
+ sky130_fd_sc_hd__dfxtp_1
X_12371_ net456 _05217_ _05226_ _05221_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__o211a_1
X_21569_ _03299_ _03300_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14110_ _06640_ _06637_ top_inst.grid_inst.data_path_wires\[3\]\[7\] VGND VGND VPWR
+ VPWR _06825_ sky130_fd_sc_hd__o21ai_4
X_23308_ net462 _04765_ _04768_ _04769_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15090_ _07733_ _07732_ VGND VGND VPWR VPWR _07740_ sky130_fd_sc_hd__nor2_1
XFILLER_0_239_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24288_ clknet_leaf_10_clk _00821_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14041_ _06735_ _06736_ _06757_ VGND VGND VPWR VPWR _06758_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_127_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23239_ net693 _04726_ _04729_ _04730_ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__o211a_1
XFILLER_0_197_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17800_ _10290_ _10291_ _10306_ VGND VGND VPWR VPWR _10308_ sky130_fd_sc_hd__and3_1
XTAP_6464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15992_ _08594_ _08565_ _08599_ VGND VGND VPWR VPWR _08601_ sky130_fd_sc_hd__nand3_1
XFILLER_0_98_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18780_ _05887_ _11205_ _11206_ _11207_ VGND VGND VPWR VPWR _11208_ sky130_fd_sc_hd__a31o_1
XTAP_6475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14943_ _07610_ _07611_ _07612_ _07092_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__o211a_1
X_17731_ _10032_ _10052_ _10050_ _10035_ VGND VGND VPWR VPWR _10240_ sky130_fd_sc_hd__a22o_1
XTAP_5774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_234_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14874_ _07546_ _07520_ VGND VGND VPWR VPWR _07558_ sky130_fd_sc_hd__and2b_1
X_17662_ _10171_ _10172_ _10032_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[2\]
+ VGND VGND VPWR VPWR _10173_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19401_ _01234_ _01235_ _01229_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__a21o_1
X_16613_ top_inst.skew_buff_inst.row\[2\].output_reg\[0\] top_inst.axis_in_inst.inbuf_bus\[16\]
+ _07059_ VGND VGND VPWR VPWR _09186_ sky130_fd_sc_hd__mux2_4
XFILLER_0_202_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13825_ _06565_ _06566_ VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__nand2_1
X_17593_ _10106_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16544_ _08876_ _08679_ _09081_ VGND VGND VPWR VPWR _09120_ sky130_fd_sc_hd__o21a_1
X_19332_ _11684_ _11679_ _11682_ _11687_ VGND VGND VPWR VPWR _11726_ sky130_fd_sc_hd__nand4_2
XFILLER_0_58_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13756_ _06455_ _06456_ VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__or2b_1
XFILLER_0_70_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12707_ _05484_ _05485_ _05516_ _05517_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_169_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16475_ _09051_ _09052_ VGND VGND VPWR VPWR _09053_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19263_ net957 _11662_ _11675_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__o21a_1
X_13687_ _06427_ _06432_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15426_ _08036_ _08035_ VGND VGND VPWR VPWR _08068_ sky130_fd_sc_hd__or2b_1
XFILLER_0_128_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18214_ _10670_ _10674_ VGND VGND VPWR VPWR _10683_ sky130_fd_sc_hd__and2b_1
X_12638_ _05447_ _05449_ _05271_ _05278_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__or4b_1
XFILLER_0_183_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19194_ _11574_ VGND VGND VPWR VPWR _11611_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15357_ _07989_ _07965_ _08000_ VGND VGND VPWR VPWR _08001_ sky130_fd_sc_hd__a21o_1
X_18145_ _10617_ _10618_ _08181_ VGND VGND VPWR VPWR _10619_ sky130_fd_sc_hd__o21ai_1
X_12569_ _05377_ _05382_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__xor2_1
XFILLER_0_182_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14308_ _07015_ _07017_ VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18076_ _05787_ _10575_ _04867_ VGND VGND VPWR VPWR _10576_ sky130_fd_sc_hd__a21oi_4
Xhold206 _00920_ VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__dlygate4sd3_1
X_15288_ _07887_ _07891_ _07889_ VGND VGND VPWR VPWR _07934_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_13_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold217 _00171_ VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 top_inst.axis_out_inst.out_buff_data\[123\] VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17027_ _09449_ _09492_ _09532_ _09576_ VGND VGND VPWR VPWR _09580_ sky130_fd_sc_hd__or4b_4
X_14239_ _06948_ _06949_ VGND VGND VPWR VPWR _06951_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold239 _00210_ VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ _11147_ _11154_ VGND VGND VPWR VPWR _11400_ sky130_fd_sc_hd__nand2_4
XFILLER_0_20_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _10418_ _10433_ VGND VGND VPWR VPWR _10434_ sky130_fd_sc_hd__xor2_1
XFILLER_0_213_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20940_ _02662_ _02708_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_205_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20871_ _02518_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__buf_4
XFILLER_0_220_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22610_ _04262_ _04265_ _04264_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__a21o_1
XFILLER_0_193_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23590_ clknet_leaf_101_clk _00123_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22541_ _04218_ _04219_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22472_ _04089_ _04153_ _04154_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24211_ clknet_leaf_17_clk _00744_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21423_ _03115_ _03116_ _03157_ _01984_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__a31o_1
XFILLER_0_228_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24142_ clknet_leaf_14_clk _00675_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21354_ top_inst.grid_inst.data_path_wires\[17\]\[2\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_241_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20305_ _02092_ _02093_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__xor2_4
X_24073_ clknet_leaf_114_clk _00606_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold740 top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[17\] VGND VGND
+ VPWR VPWR net922 sky130_fd_sc_hd__dlygate4sd3_1
X_21285_ _02993_ _02994_ _03022_ _03023_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__a211o_1
XFILLER_0_188_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold751 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[20\] VGND
+ VGND VPWR VPWR net933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold762 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[28\] VGND
+ VGND VPWR VPWR net944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23024_ net951 _04603_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold773 top_inst.axis_out_inst.out_buff_data\[15\] VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__dlygate4sd3_1
X_20236_ _01990_ _01987_ _02009_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__and3_1
XFILLER_0_229_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold784 top_inst.deskew_buff_inst.col_input\[51\] VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold795 top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[1\] VGND VGND
+ VPWR VPWR net977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_244_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20167_ _01950_ _01958_ _01976_ _01939_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__a22o_1
XFILLER_0_244_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20098_ _01884_ _01864_ _01906_ _01910_ _01905_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__a32o_1
XTAP_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23926_ clknet_leaf_76_clk _00459_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ net610 _04969_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__or2_1
XFILLER_0_207_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_212_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23857_ clknet_leaf_68_clk _00390_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[13\] _04930_
+ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__or2_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _06355_ _06357_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__xnor2_1
X_22808_ _04464_ _04475_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__xnor2_1
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _07278_ _07280_ VGND VGND VPWR VPWR _07281_ sky130_fd_sc_hd__nor2_4
XFILLER_0_79_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23788_ clknet_leaf_70_clk _00321_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13541_ _06272_ _06275_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__nand2_1
X_22739_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[25\] _04215_ _04216_
+ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_67_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16260_ _08841_ _08842_ VGND VGND VPWR VPWR _08843_ sky130_fd_sc_hd__nand2_1
X_13472_ _06223_ _06224_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15211_ _07805_ _07807_ VGND VGND VPWR VPWR _07859_ sky130_fd_sc_hd__and2b_1
XFILLER_0_124_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24409_ clknet_leaf_57_clk _00942_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12423_ net288 _05243_ _05255_ _05247_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16191_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[5\] _08775_ VGND
+ VGND VPWR VPWR _08776_ sky130_fd_sc_hd__xor2_2
XFILLER_0_30_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15142_ _07789_ _07790_ VGND VGND VPWR VPWR _07791_ sky130_fd_sc_hd__nand2_1
X_12354_ net691 _05204_ _05216_ _05208_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_244_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19950_ _01611_ _01743_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__nor2_2
X_15073_ _07722_ _07723_ VGND VGND VPWR VPWR _07724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12285_ _04858_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__clkbuf_8
X_14024_ _06652_ _06650_ _06622_ top_inst.grid_inst.data_path_wires\[3\]\[0\] VGND
+ VGND VPWR VPWR _06741_ sky130_fd_sc_hd__nand4_4
X_18901_ _11284_ _11286_ VGND VGND VPWR VPWR _11325_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19881_ _01697_ _01703_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__xnor2_2
X_18832_ _11257_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__clkbuf_1
XTAP_6250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1032 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_234_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18763_ _11182_ _11183_ VGND VGND VPWR VPWR _11191_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15975_ _08582_ _08584_ VGND VGND VPWR VPWR _08585_ sky130_fd_sc_hd__nand2_1
XTAP_5571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17714_ _10184_ _10223_ VGND VGND VPWR VPWR _10224_ sky130_fd_sc_hd__xor2_1
X_14926_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[24\] _07576_ VGND
+ VGND VPWR VPWR _07602_ sky130_fd_sc_hd__and2_1
XFILLER_0_175_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18694_ top_inst.grid_inst.data_path_wires\[13\]\[3\] VGND VGND VPWR VPWR _11138_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_117_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17645_ _10139_ _10135_ VGND VGND VPWR VPWR _10156_ sky130_fd_sc_hd__or2b_1
X_14857_ _07540_ _07541_ VGND VGND VPWR VPWR _07542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_203_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_216_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13808_ _06522_ _06519_ _06550_ VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__a21o_1
X_14788_ _07448_ _07473_ _07474_ VGND VGND VPWR VPWR _07475_ sky130_fd_sc_hd__and3_1
X_17576_ _10087_ _10089_ VGND VGND VPWR VPWR _10090_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19315_ _11679_ _11677_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _11711_ sky130_fd_sc_hd__a21oi_1
X_16527_ _09054_ _09059_ _09057_ VGND VGND VPWR VPWR _09104_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13739_ _06483_ VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19246_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[16\] _10639_ VGND
+ VGND VPWR VPWR _11661_ sky130_fd_sc_hd__or2_1
X_16458_ _09035_ _09036_ VGND VGND VPWR VPWR _09037_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15409_ _08003_ _08010_ _08001_ VGND VGND VPWR VPWR _08052_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_171_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16389_ _08677_ _08967_ _08968_ VGND VGND VPWR VPWR _08969_ sky130_fd_sc_hd__a21bo_1
X_19177_ _11589_ _11593_ VGND VGND VPWR VPWR _11594_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18128_ top_inst.grid_inst.data_path_wires\[12\]\[4\] VGND VGND VPWR VPWR _10606_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18059_ _10536_ _10559_ VGND VGND VPWR VPWR _10560_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_223_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21070_ _02832_ _02833_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__xor2_1
XFILLER_0_223_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20021_ _01824_ _01837_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__xor2_2
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21972_ _02864_ _02877_ _03683_ _03660_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer10 net190 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_1
Xrebuffer21 _09214_ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__buf_6
XFILLER_0_154_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer32 _09522_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23711_ clknet_leaf_124_clk _00244_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_234_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20923_ _02645_ _02692_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer43 net224 VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer54 _01282_ VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer65 net246 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_16_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer76 net1122 VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__clkbuf_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23642_ clknet_leaf_127_clk _00175_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20854_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[18\] _02559_ _02600_
+ _02598_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23573_ clknet_leaf_129_clk _00106_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20785_ _02558_ _02560_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22524_ _04189_ _04190_ _04204_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_130_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22455_ _04135_ _04100_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21406_ top_inst.grid_inst.data_path_wires\[17\]\[2\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[6\]
+ _03090_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22386_ _04067_ _04070_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_241_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24125_ clknet_leaf_119_clk _00658_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_114_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21337_ _03036_ _03042_ _03073_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24056_ clknet_leaf_46_clk _00589_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_12070_ net481 _05050_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__or2_1
Xhold570 top_inst.axis_out_inst.out_buff_data\[60\] VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__dlygate4sd3_1
X_21268_ _02965_ _02970_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__or2b_1
XFILLER_0_241_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold581 top_inst.axis_out_inst.out_buff_data\[45\] VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold592 top_inst.axis_out_inst.out_buff_data\[18\] VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__dlygate4sd3_1
X_23007_ net1019 _04588_ _04595_ _04590_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__o211a_1
X_20219_ _02015_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21199_ top_inst.deskew_buff_inst.col_input\[67\] _05730_ VGND VGND VPWR VPWR _02941_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_217_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_216_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_232_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[8\] _08374_ VGND
+ VGND VPWR VPWR _08375_ sky130_fd_sc_hd__xnor2_1
X_12972_ _05763_ _05294_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__or2_1
XTAP_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _07398_ _07399_ VGND VGND VPWR VPWR _07400_ sky130_fd_sc_hd__and2_1
XTAP_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11923_ top_inst.axis_out_inst.out_buff_data\[35\] _04969_ VGND VGND VPWR VPWR _04971_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_73_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23909_ clknet_leaf_36_clk _00442_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15691_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[6\] _08306_ _08307_
+ VGND VGND VPWR VPWR _08308_ sky130_fd_sc_hd__mux2_1
XTAP_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14642_ _07328_ _07331_ VGND VGND VPWR VPWR _07332_ sky130_fd_sc_hd__xor2_1
X_17430_ _09951_ _09967_ VGND VGND VPWR VPWR _09968_ sky130_fd_sc_hd__xnor2_1
XTAP_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ net362 _04930_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__or2_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17361_ _09893_ _09901_ VGND VGND VPWR VPWR _09902_ sky130_fd_sc_hd__xnor2_2
X_14573_ _07217_ _07263_ _07264_ VGND VGND VPWR VPWR _07265_ sky130_fd_sc_hd__and3_1
XFILLER_0_185_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11785_ net337 _04885_ _04892_ _04889_ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19100_ _11512_ _11518_ VGND VGND VPWR VPWR _11519_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16312_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[1\] _08682_ top_inst.grid_inst.data_path_wires\[8\]\[7\]
+ VGND VGND VPWR VPWR _08894_ sky130_fd_sc_hd__o21ai_2
X_13524_ top_inst.grid_inst.data_path_wires\[2\]\[4\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[2\]\[5\]
+ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__a22oi_1
X_17292_ _09623_ _09835_ VGND VGND VPWR VPWR _09836_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16243_ _08736_ _08758_ _08783_ _08787_ VGND VGND VPWR VPWR _08827_ sky130_fd_sc_hd__o31a_1
X_19031_ _11450_ _11451_ VGND VGND VPWR VPWR _11452_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13455_ _06212_ _05773_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12406_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[19\] _05235_
+ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__or2_1
X_16174_ _08758_ _08759_ VGND VGND VPWR VPWR _08760_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13386_ _06113_ _06158_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15125_ _07773_ _07774_ VGND VGND VPWR VPWR _07775_ sky130_fd_sc_hd__nor2_1
Xoutput108 net108 VGND VGND VPWR VPWR output_tdata[48] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12337_ net298 _05196_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__or2_1
Xoutput119 net119 VGND VGND VPWR VPWR output_tdata[58] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15056_ _07707_ VGND VGND VPWR VPWR _07708_ sky130_fd_sc_hd__clkbuf_8
X_19933_ _01652_ _01751_ _01753_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__a21o_1
XFILLER_0_220_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12268_ _05127_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__buf_2
XFILLER_0_208_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_1296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14007_ _06670_ _06686_ _06687_ _06724_ VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__a31o_1
X_19864_ _01682_ _01687_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__xor2_2
XFILLER_0_120_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12199_ net526 _05123_ _05126_ _05128_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__o211a_1
Xoutput90 net90 VGND VGND VPWR VPWR output_tdata[31] sky130_fd_sc_hd__clkbuf_4
X_18815_ top_inst.grid_inst.data_path_wires\[13\]\[5\] top_inst.grid_inst.data_path_wires\[13\]\[4\]
+ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _11241_ sky130_fd_sc_hd__nand4_1
XFILLER_0_235_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19795_ _01594_ _01595_ _01621_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_170_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18746_ _11174_ _11175_ _06682_ VGND VGND VPWR VPWR _11176_ sky130_fd_sc_hd__a21o_1
XTAP_5390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15958_ _08557_ _08525_ _08567_ VGND VGND VPWR VPWR _08568_ sky130_fd_sc_hd__a21o_1
X_14909_ _07578_ _07590_ _07591_ _05315_ VGND VGND VPWR VPWR _07592_ sky130_fd_sc_hd__and4b_2
XFILLER_0_37_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18677_ net1046 _11116_ net167 VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15889_ _08499_ _08500_ VGND VGND VPWR VPWR _08501_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_231_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17628_ _10135_ _10139_ VGND VGND VPWR VPWR _10140_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_1272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17559_ _10027_ _10025_ _10044_ _10042_ VGND VGND VPWR VPWR _10074_ sky130_fd_sc_hd__nand4_1
XFILLER_0_58_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_1346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20570_ _02312_ _02341_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19229_ _11479_ VGND VGND VPWR VPWR _11644_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22240_ _02706_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__buf_4
XFILLER_0_108_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1015 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22171_ top_inst.grid_inst.data_path_wires\[18\]\[4\] _03705_ _03686_ _03707_ VGND
+ VGND VPWR VPWR _03861_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21122_ _02001_ _11142_ _02876_ _02707_ VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21053_ _02816_ _02817_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20004_ _01788_ net168 VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1014 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21955_ _03665_ _03652_ _03668_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__a21o_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20906_ _02673_ _02676_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__xnor2_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1057 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21886_ _03603_ _03604_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_234_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23625_ clknet_leaf_102_clk net265 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20837_ _02586_ _02610_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__xor2_1
XFILLER_0_132_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23556_ clknet_leaf_102_clk _00089_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20768_ net270 _01386_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22507_ _04053_ _04185_ _04186_ _04187_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23487_ clknet_leaf_141_clk _00020_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[77\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20699_ _02437_ _02441_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__and2b_1
XFILLER_0_208_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13240_ _05750_ _05765_ _05763_ top_inst.grid_inst.data_path_wires\[1\]\[7\] VGND
+ VGND VPWR VPWR _06017_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_134_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22438_ _04091_ _04121_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__xor2_1
XFILLER_0_123_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13171_ _05944_ _05906_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22369_ _04042_ _04044_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24108_ clknet_leaf_14_clk _00641_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_12122_ _05044_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_104_1414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1059 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16930_ _09483_ _09484_ _09439_ _09458_ VGND VGND VPWR VPWR _09486_ sky130_fd_sc_hd__o211ai_1
X_24039_ clknet_leaf_42_clk _00572_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_12053_ _05044_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16861_ _09193_ _09188_ net219 VGND VGND VPWR VPWR _09418_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_232_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18600_ _11058_ _11059_ VGND VGND VPWR VPWR _11060_ sky130_fd_sc_hd__nor2_1
XFILLER_0_189_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15812_ _08424_ _08425_ VGND VGND VPWR VPWR _08426_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_217_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19580_ _01363_ _01365_ _01364_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_137_1212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16792_ _09348_ _09349_ net170 _09316_ VGND VGND VPWR VPWR _09351_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_232_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18531_ _10991_ _10992_ VGND VGND VPWR VPWR _10993_ sky130_fd_sc_hd__nand2_1
X_12955_ _05739_ _05641_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__nand2_1
X_15743_ _08313_ _08314_ VGND VGND VPWR VPWR _08358_ sky130_fd_sc_hd__nor2_1
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[28\] _04956_
+ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__or2_1
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18462_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[11\] _10793_ VGND
+ VGND VPWR VPWR _10925_ sky130_fd_sc_hd__xnor2_1
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _05660_ _05670_ _05690_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__nand3_1
XFILLER_0_59_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _08289_ _08290_ VGND VGND VPWR VPWR _08291_ sky130_fd_sc_hd__and2_1
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _09942_ _09943_ VGND VGND VPWR VPWR _09951_ sky130_fd_sc_hd__or2b_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14625_ _07306_ _07307_ VGND VGND VPWR VPWR _07315_ sky130_fd_sc_hd__and2b_1
XFILLER_0_184_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11837_ top_inst.axis_out_inst.out_buff_data\[94\] _04917_ VGND VGND VPWR VPWR _04922_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_96_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_213_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18393_ top_inst.grid_inst.data_path_wires\[12\]\[3\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[6\]
+ _10857_ top_inst.grid_inst.data_path_wires\[12\]\[2\] VGND VGND VPWR VPWR _10858_
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _07245_ _07246_ _07205_ VGND VGND VPWR VPWR _07248_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17344_ _07707_ VGND VGND VPWR VPWR _09886_ sky130_fd_sc_hd__clkbuf_8
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ net625 _04860_ _04882_ _04875_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_891 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13507_ _06235_ _06257_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__xor2_1
X_17275_ _09808_ _09818_ _09810_ VGND VGND VPWR VPWR _09820_ sky130_fd_sc_hd__nand3_1
X_14487_ _07178_ _07179_ net1125 VGND VGND VPWR VPWR _07181_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_181_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_859 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19014_ _11431_ _11434_ VGND VGND VPWR VPWR _11435_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16226_ _08676_ top_inst.grid_inst.data_path_wires\[8\]\[5\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[1\]
+ _08682_ VGND VGND VPWR VPWR _08810_ sky130_fd_sc_hd__nand4_1
X_13438_ _06200_ _05773_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__or2_1
Xrebuffer1 _09446_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__buf_1
XFILLER_0_140_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16157_ top_inst.grid_inst.data_path_wires\[8\]\[3\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[1\]
+ _08682_ top_inst.grid_inst.data_path_wires\[8\]\[4\] VGND VGND VPWR VPWR _08743_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13369_ _06139_ _06142_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[13\]
+ _05327_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_12_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15108_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[6\] _07756_ _07757_
+ VGND VGND VPWR VPWR _07758_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16088_ _08661_ _08681_ _08685_ _08666_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19916_ _01721_ _01724_ _01723_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__a21o_1
X_15039_ _07689_ _07690_ VGND VGND VPWR VPWR _07691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19847_ _01642_ _01670_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_235_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1000 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_1155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19778_ _01298_ _11709_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18729_ _11143_ _10607_ _11162_ _11160_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21740_ net878 _02491_ _03464_ _03465_ _02962_ VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__o221a_1
XFILLER_0_17_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21671_ _03394_ _03399_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23410_ net530 _04655_ _04825_ _04819_ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20622_ _02395_ _02402_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__xor2_1
X_24390_ clknet_leaf_38_clk _00923_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_1007 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23341_ net619 _04778_ _04787_ _04782_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20553_ _02334_ _02335_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__xor2_1
XFILLER_0_117_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23272_ net364 _04739_ _04748_ _04743_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20484_ _02267_ _02264_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22223_ _03823_ _03870_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_972 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22154_ top_inst.deskew_buff_inst.col_input\[102\] _03844_ _06140_ VGND VGND VPWR
+ VPWR _03845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21105_ _02864_ _11133_ VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__or2_1
X_22085_ _03753_ _03773_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_196_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_1__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_4_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_21036_ _02763_ _02783_ _02801_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_1407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22987_ net902 _04575_ _04584_ _04577_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12740_ _05545_ _05549_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__and2_2
XFILLER_0_215_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21938_ _03652_ _03653_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _05482_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21869_ _03587_ _03588_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__nor2_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _07105_ _07106_ VGND VGND VPWR VPWR _07107_ sky130_fd_sc_hd__nand2_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23608_ clknet_leaf_103_clk net459 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15390_ _07622_ _07824_ _08031_ VGND VGND VPWR VPWR _08033_ sky130_fd_sc_hd__nor3_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24588_ clknet_leaf_32_clk _01121_ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_65_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14341_ _07043_ _07044_ _07041_ VGND VGND VPWR VPWR _07049_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23539_ clknet_leaf_131_clk _00072_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17060_ _09611_ _09612_ VGND VGND VPWR VPWR _09613_ sky130_fd_sc_hd__xnor2_2
X_14272_ _06943_ _06947_ _06941_ VGND VGND VPWR VPWR _06983_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16011_ _08618_ _08619_ VGND VGND VPWR VPWR _08620_ sky130_fd_sc_hd__nor2_2
XFILLER_0_180_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13223_ _05998_ _06000_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13154_ _05889_ _05890_ _05932_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_20_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _04994_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_130_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ top_inst.grid_inst.data_path_wires\[1\]\[5\] _05759_ _05757_ _05750_ VGND
+ VGND VPWR VPWR _05866_ sky130_fd_sc_hd__a22oi_1
X_17962_ _10464_ _10465_ VGND VGND VPWR VPWR _10466_ sky130_fd_sc_hd__and2_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19701_ _01528_ _01529_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__xor2_1
X_16913_ _09465_ _09468_ VGND VGND VPWR VPWR _09469_ sky130_fd_sc_hd__xor2_1
X_12036_ net966 _05031_ _05034_ _05035_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__o211a_1
XFILLER_0_224_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17893_ _10397_ _10398_ VGND VGND VPWR VPWR _10399_ sky130_fd_sc_hd__and2_1
XFILLER_0_217_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19632_ _01460_ _01461_ _01434_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__a21oi_1
X_16844_ _09398_ _09400_ _09350_ VGND VGND VPWR VPWR _09402_ sky130_fd_sc_hd__a21o_1
XFILLER_0_233_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19563_ _01394_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__buf_2
X_16775_ _09207_ _09203_ _09197_ _09202_ VGND VGND VPWR VPWR _09334_ sky130_fd_sc_hd__nand4_2
XFILLER_0_87_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13987_ _06676_ _06696_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18514_ _10589_ _10857_ VGND VGND VPWR VPWR _10976_ sky130_fd_sc_hd__nor2_1
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15726_ _08300_ _08341_ VGND VGND VPWR VPWR _08342_ sky130_fd_sc_hd__xor2_1
X_12938_ _05739_ _05488_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__nand2_1
X_19494_ _01325_ _01326_ _01327_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18445_ _10907_ _10908_ VGND VGND VPWR VPWR _10909_ sky130_fd_sc_hd__xnor2_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15657_ top_inst.grid_inst.data_path_wires\[7\]\[0\] _08169_ _08167_ _08137_ VGND
+ VGND VPWR VPWR _08274_ sky130_fd_sc_hd__a22o_1
X_12869_ _05673_ _05674_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__or2_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14608_ _07289_ _07298_ VGND VGND VPWR VPWR _07299_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18376_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[8\] _10793_ _10840_
+ VGND VGND VPWR VPWR _10841_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15588_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[2\] _08184_ _08185_
+ VGND VGND VPWR VPWR _08208_ sky130_fd_sc_hd__a21boi_2
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17327_ _09726_ _09855_ VGND VGND VPWR VPWR _09869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14539_ _07066_ _07229_ _07230_ VGND VGND VPWR VPWR _07231_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_43_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17258_ _06701_ VGND VGND VPWR VPWR _09804_ sky130_fd_sc_hd__buf_4
XFILLER_0_153_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16209_ _08780_ _08782_ VGND VGND VPWR VPWR _08793_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17189_ _09727_ _09737_ VGND VGND VPWR VPWR _09738_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_236_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22910_ net766 _04535_ _04540_ _04537_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23890_ clknet_leaf_62_clk _00423_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22841_ net898 _04496_ _04501_ _04498_ VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22772_ _04409_ _04421_ _04441_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24511_ clknet_leaf_132_clk _01044_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dfxtp_4
X_21723_ _03278_ _03448_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_231_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24442_ clknet_leaf_64_clk net984 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[0\].output_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21654_ _03375_ _03382_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20605_ _02262_ _02308_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__or2_1
X_24373_ clknet_leaf_38_clk net899 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].output_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21585_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[14\] _03080_ VGND
+ VGND VPWR VPWR _03316_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_954 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23324_ net415 _04765_ _04777_ _04769_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20536_ _01995_ _02229_ _02317_ _02318_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__o22a_1
XFILLER_0_127_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23255_ net920 _04726_ _04738_ _04730_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20467_ _02248_ _02249_ _02250_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22206_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[8\] _03894_ VGND
+ VGND VPWR VPWR _03895_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23186_ net736 _04685_ _04699_ _04691_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20398_ _02177_ _02183_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__xnor2_1
XTAP_6602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22137_ _03688_ _03703_ _03825_ _03826_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__o2bb2a_1
XTAP_6624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22068_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[4\] _03760_ VGND
+ VGND VPWR VPWR _03761_ sky130_fd_sc_hd__xor2_2
XTAP_6679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13910_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[1\] VGND VGND
+ VPWR VPWR _06640_ sky130_fd_sc_hd__clkbuf_4
X_21019_ _02643_ _02766_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__and2_1
XTAP_5978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14890_ _07557_ _07573_ VGND VGND VPWR VPWR _07574_ sky130_fd_sc_hd__nor2_1
XTAP_5989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1063 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13841_ _06140_ _06582_ VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__nand2_1
XFILLER_0_230_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16560_ _09093_ _09097_ _09095_ VGND VGND VPWR VPWR _09136_ sky130_fd_sc_hd__a21oi_2
X_13772_ _06470_ _06472_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15511_ _08145_ _04859_ VGND VGND VPWR VPWR _08146_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12723_ _05492_ _05493_ _05491_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16491_ _09066_ _09068_ VGND VGND VPWR VPWR _09069_ sky130_fd_sc_hd__and2_1
XFILLER_0_195_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18230_ _10690_ _10698_ VGND VGND VPWR VPWR _10699_ sky130_fd_sc_hd__xor2_2
X_12654_ _05304_ _05463_ _05465_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__and3_1
X_15442_ _08067_ _08049_ _08083_ VGND VGND VPWR VPWR _08084_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_242_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18161_ _10622_ _10623_ VGND VGND VPWR VPWR _10633_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15373_ _07978_ _07980_ VGND VGND VPWR VPWR _08017_ sky130_fd_sc_hd__or2b_1
X_12585_ _05325_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__buf_8
XFILLER_0_53_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17112_ _09622_ _09616_ _09657_ VGND VGND VPWR VPWR _09663_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14324_ _07002_ _07005_ _07031_ VGND VGND VPWR VPWR _07033_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18092_ _10025_ _08663_ _10580_ _10448_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17043_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[5\] net219 VGND
+ VGND VPWR VPWR _09596_ sky130_fd_sc_hd__and2_1
X_14255_ _06635_ _06650_ VGND VGND VPWR VPWR _06966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13206_ _05937_ _05938_ _05934_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__or3b_1
XFILLER_0_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_1268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14186_ top_inst.grid_inst.data_path_wires\[3\]\[6\] _06648_ _06645_ _06635_ VGND
+ VGND VPWR VPWR _06899_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13137_ _05872_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__inv_2
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18994_ _11413_ _11415_ VGND VGND VPWR VPWR _11416_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _05831_ _05834_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__nand2_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _10397_ _10439_ _10440_ VGND VGND VPWR VPWR _10449_ sky130_fd_sc_hd__or3_1
XFILLER_0_104_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12019_ net439 _05023_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__or2_1
XFILLER_0_224_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17876_ _10380_ VGND VGND VPWR VPWR _10382_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19615_ _01297_ _01314_ _11691_ _11695_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__or4b_4
X_16827_ _09382_ _09383_ _09375_ VGND VGND VPWR VPWR _09385_ sky130_fd_sc_hd__a21o_1
XFILLER_0_233_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19546_ _01376_ _01377_ _01323_ _01325_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16758_ _09316_ _09317_ VGND VGND VPWR VPWR _09318_ sky130_fd_sc_hd__or2_4
XFILLER_0_220_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15709_ _08149_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[1\] _08154_
+ top_inst.grid_inst.data_path_wires\[7\]\[7\] VGND VGND VPWR VPWR _08325_ sky130_fd_sc_hd__a22o_1
X_19477_ _01309_ _01310_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__nor2_1
XFILLER_0_220_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16689_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[3\] _09250_ VGND
+ VGND VPWR VPWR _09251_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18428_ top_inst.grid_inst.data_path_wires\[12\]\[7\] _10608_ _10604_ VGND VGND VPWR
+ VPWR _10892_ sky130_fd_sc_hd__and3_1
XFILLER_0_173_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18359_ _10822_ _10824_ VGND VGND VPWR VPWR _10825_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21370_ _03059_ _03034_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20321_ top_inst.grid_inst.data_path_wires\[16\]\[4\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[1\]
+ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold900 top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[17\] VGND VGND
+ VPWR VPWR net1082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 top_inst.deskew_buff_inst.col_input\[15\] VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold922 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[11\] VGND
+ VGND VPWR VPWR net1104 sky130_fd_sc_hd__dlygate4sd3_1
X_23040_ _04600_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold933 top_inst.axis_in_inst.inbuf_bus\[30\] VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__dlygate4sd3_1
X_20252_ _02029_ _02042_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__xor2_1
XFILLER_0_228_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20183_ _10030_ _11682_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__or2_1
XFILLER_0_228_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23942_ clknet_leaf_81_clk _00475_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_1203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23873_ clknet_leaf_50_clk _00406_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22824_ _04092_ _04268_ _04489_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[27\]
+ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__a31o_1
XFILLER_0_233_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22755_ _04417_ _04418_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__or2b_1
XFILLER_0_165_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xsplit37 _09218_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21706_ _03431_ _03432_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22686_ net608 _03528_ _04358_ _04359_ _09806_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__o221a_1
XFILLER_0_168_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24425_ clknet_leaf_57_clk net735 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].output_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21637_ _03347_ _03343_ _03366_ VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24356_ clknet_leaf_26_clk _00889_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[115\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12370_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[3\] _05222_
+ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21568_ _03249_ _03250_ _03264_ _03263_ _03261_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__o32a_1
XFILLER_0_145_691 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23307_ _04690_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20519_ _02271_ _02301_ _02302_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__and3_1
X_24287_ clknet_leaf_10_clk _00820_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_166_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21499_ _03197_ _03193_ _03231_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14040_ _06738_ _06756_ VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__xor2_1
XFILLER_0_160_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23238_ _04690_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_240_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23169_ _04690_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__clkbuf_4
XTAP_6421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ _08594_ _08565_ _08599_ VGND VGND VPWR VPWR _08600_ sky130_fd_sc_hd__a21oi_1
XTAP_6476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17730_ _10232_ _10238_ VGND VGND VPWR VPWR _10239_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14942_ _05739_ _07290_ VGND VGND VPWR VPWR _07612_ sky130_fd_sc_hd__nand2_1
XTAP_5764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17661_ top_inst.grid_inst.data_path_wires\[11\]\[3\] top_inst.grid_inst.data_path_wires\[11\]\[2\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _10172_ sky130_fd_sc_hd__and4_1
XFILLER_0_215_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14873_ _07550_ _07552_ _07556_ VGND VGND VPWR VPWR _07557_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_202_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19400_ _01229_ _01234_ _01235_ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__nand3_2
XFILLER_0_72_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16612_ _05269_ VGND VGND VPWR VPWR _09185_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_203_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13824_ _06496_ _06564_ VGND VGND VPWR VPWR _06566_ sky130_fd_sc_hd__or2_1
XFILLER_0_230_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17592_ _09661_ _10105_ VGND VGND VPWR VPWR _10106_ sky130_fd_sc_hd__and2_1
XFILLER_0_202_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19331_ _11684_ _11682_ _11687_ _11679_ VGND VGND VPWR VPWR _11725_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16543_ _09040_ _09082_ _09083_ VGND VGND VPWR VPWR _09119_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_70_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_202_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13755_ _06497_ _06498_ VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12706_ _05486_ _05487_ _05515_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__and3_1
XFILLER_0_183_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19262_ net963 _11662_ _11675_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__o21a_1
X_16474_ _09039_ _09015_ _09050_ VGND VGND VPWR VPWR _09052_ sky130_fd_sc_hd__nand3_1
XFILLER_0_195_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_956 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13686_ _06430_ _06431_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18213_ _10659_ _10678_ VGND VGND VPWR VPWR _10682_ sky130_fd_sc_hd__nor2_1
X_15425_ _08030_ _07998_ _08040_ VGND VGND VPWR VPWR _08067_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12637_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _05449_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19193_ _11587_ _11609_ VGND VGND VPWR VPWR _11610_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18144_ _10577_ _10597_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _10618_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12568_ _05380_ _05381_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__xor2_1
XFILLER_0_142_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15356_ _07998_ _07999_ VGND VGND VPWR VPWR _08000_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_842 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14307_ _06945_ _06984_ _07016_ VGND VGND VPWR VPWR _07017_ sky130_fd_sc_hd__a21oi_1
X_18075_ _10544_ _10560_ _10573_ _10574_ VGND VGND VPWR VPWR _10575_ sky130_fd_sc_hd__a211o_1
X_12499_ _05273_ _05272_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15287_ _07930_ _07932_ VGND VGND VPWR VPWR _07933_ sky130_fd_sc_hd__xnor2_2
Xhold207 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[5\] VGND VGND
+ VPWR VPWR net389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold218 top_inst.deskew_buff_inst.col_input\[30\] VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__buf_1
X_17026_ _09532_ _09576_ VGND VGND VPWR VPWR _09579_ sky130_fd_sc_hd__or2b_1
Xhold229 top_inst.deskew_buff_inst.col_input\[80\] VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ _06948_ _06949_ VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14169_ _06881_ _06882_ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__or2b_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _11396_ _11398_ VGND VGND VPWR VPWR _11399_ sky130_fd_sc_hd__and2_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _10430_ _10432_ VGND VGND VPWR VPWR _10433_ sky130_fd_sc_hd__xor2_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17859_ _10330_ _10329_ VGND VGND VPWR VPWR _10365_ sky130_fd_sc_hd__or2b_1
XFILLER_0_234_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20870_ _02626_ _02627_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19529_ _01358_ _01361_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22540_ _04218_ _04219_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22471_ _04083_ _04090_ _04120_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_228_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24210_ clknet_leaf_17_clk _00743_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21422_ _03115_ _03116_ _03157_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_161_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24141_ clknet_leaf_144_clk _00674_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21353_ top_inst.grid_inst.data_path_wires\[17\]\[1\] _02897_ VGND VGND VPWR VPWR
+ _03090_ sky130_fd_sc_hd__and2b_1
XFILLER_0_163_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20304_ _02062_ _02063_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__nor2b_2
X_24072_ clknet_leaf_114_clk _00605_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold730 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[4\] VGND
+ VGND VPWR VPWR net912 sky130_fd_sc_hd__dlygate4sd3_1
X_21284_ _03020_ _03021_ _02995_ _02996_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__o211a_1
Xhold741 top_inst.deskew_buff_inst.col_input\[113\] VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23023_ net12 _04601_ _04605_ _04606_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__o211a_1
Xhold752 top_inst.deskew_buff_inst.col_input\[23\] VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold763 top_inst.axis_out_inst.out_buff_data\[55\] VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__dlygate4sd3_1
X_20235_ _01987_ _02009_ _02007_ _01990_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__a22o_1
Xhold774 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[18\] VGND VGND
+ VPWR VPWR net956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold785 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[16\] VGND
+ VGND VPWR VPWR net967 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold796 top_inst.axis_out_inst.out_buff_data\[52\] VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20166_ _01783_ _01956_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20097_ _01879_ _01882_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__nand2_1
XTAP_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23925_ clknet_leaf_76_clk _00458_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_207_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11870_ net839 _04938_ _04940_ _04929_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__o211a_1
X_23856_ clknet_leaf_69_clk _00389_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22807_ _04466_ _04474_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23787_ clknet_leaf_70_clk _00320_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_20999_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[25\] _02666_ _02765_
+ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__o21a_1
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13540_ _06281_ _06283_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__or2_1
XFILLER_0_223_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22738_ _04364_ _04407_ _04408_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13471_ _06184_ _06202_ _06217_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__and3_1
XFILLER_0_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22669_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[21\] _04215_ _04216_
+ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__a21o_1
X_15210_ _07856_ _07857_ VGND VGND VPWR VPWR _07858_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12422_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[26\] _05248_
+ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__or2_1
X_24408_ clknet_leaf_39_clk net713 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].output_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16190_ _08773_ _08774_ VGND VGND VPWR VPWR _08775_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15141_ _07619_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[2\] _07787_
+ _07788_ VGND VGND VPWR VPWR _07790_ sky130_fd_sc_hd__nand4_2
XFILLER_0_51_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12353_ net680 _05209_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24339_ clknet_leaf_9_clk _00872_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[98\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15072_ top_inst.grid_inst.data_path_wires\[6\]\[5\] top_inst.grid_inst.data_path_wires\[6\]\[4\]
+ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[1\] _07626_ VGND VGND
+ VPWR VPWR _07723_ sky130_fd_sc_hd__nand4_1
X_12284_ net400 _05164_ _05176_ _05168_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14023_ _06650_ _06622_ _06618_ _06652_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__a22o_1
X_18900_ _11298_ _11323_ VGND VGND VPWR VPWR _11324_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19880_ _01701_ _01702_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_222_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18831_ _10641_ _11256_ VGND VGND VPWR VPWR _11257_ sky130_fd_sc_hd__and2_1
XTAP_6240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18762_ _11175_ _11187_ VGND VGND VPWR VPWR _11190_ sky130_fd_sc_hd__and2b_1
XTAP_6295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15974_ _08538_ _08539_ _08583_ VGND VGND VPWR VPWR _08584_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_234_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17713_ _10059_ _10222_ VGND VGND VPWR VPWR _10223_ sky130_fd_sc_hd__xnor2_1
X_14925_ _07593_ _07601_ _07594_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__o21a_1
XTAP_5583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18693_ _10581_ _10584_ _11136_ _11137_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__o211a_1
XFILLER_0_234_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold90 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[13\] VGND
+ VGND VPWR VPWR net272 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17644_ _10143_ _10145_ VGND VGND VPWR VPWR _10155_ sky130_fd_sc_hd__nand2_1
X_14856_ _07538_ _07539_ VGND VGND VPWR VPWR _07541_ sky130_fd_sc_hd__nand2_1
XTAP_4893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13807_ _06548_ _06549_ VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__nand2_1
X_17575_ _10047_ _10088_ VGND VGND VPWR VPWR _10089_ sky130_fd_sc_hd__nand2_2
XFILLER_0_216_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14787_ _07471_ _07472_ _07425_ _07428_ VGND VGND VPWR VPWR _07474_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_212_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11999_ net758 _05004_ _05014_ _05008_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19314_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[7\] _05276_ _11710_
+ _11641_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16526_ _09101_ _09102_ VGND VGND VPWR VPWR _09103_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13738_ _06364_ _06482_ VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19245_ _11643_ _11659_ VGND VGND VPWR VPWR _11660_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16457_ _08992_ _08994_ _08990_ VGND VGND VPWR VPWR _09036_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13669_ _06413_ _06414_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15408_ _08049_ _08050_ VGND VGND VPWR VPWR _08051_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19176_ _11514_ _11592_ VGND VGND VPWR VPWR _11593_ sky130_fd_sc_hd__xor2_1
X_16388_ _08676_ _08693_ _08690_ top_inst.grid_inst.data_path_wires\[8\]\[7\] VGND
+ VGND VPWR VPWR _08968_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18127_ _10585_ _10046_ _10605_ _10594_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__o211a_1
X_15339_ _07982_ _07983_ VGND VGND VPWR VPWR _07984_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18058_ _10556_ _10558_ VGND VGND VPWR VPWR _10559_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17009_ net1117 _09561_ _09553_ VGND VGND VPWR VPWR _09563_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_22_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20020_ _01813_ _01836_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__xor2_2
XFILLER_0_158_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21971_ _03682_ _02869_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__or2_1
XFILLER_0_213_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer11 _11699_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_6
XFILLER_0_94_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer22 _09518_ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_2
X_20922_ _02690_ _02691_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__nor2_1
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23710_ clknet_leaf_123_clk _00243_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer33 _09205_ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_1
Xrebuffer44 _09517_ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__buf_1
XFILLER_0_174_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_234_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer55 _01285_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_867 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer66 net247 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer77 _07437_ VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20853_ _02624_ _02625_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__and2_1
X_23641_ clknet_leaf_125_clk net419 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_234_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23572_ clknet_leaf_108_clk _00105_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20784_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[15\] _02559_ _02524_
+ _02522_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1027 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22523_ _04191_ _04203_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22454_ _04025_ _04136_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__nor2_4
XFILLER_0_31_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21405_ _03137_ _03140_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_161_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22385_ _04068_ _04069_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24124_ clknet_leaf_118_clk _00657_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_241_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21336_ _03037_ _03041_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__nor2_1
XFILLER_0_206_1344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1011 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24055_ clknet_leaf_34_clk _00588_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[31\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold560 top_inst.axis_out_inst.out_buff_data\[83\] VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__dlygate4sd3_1
X_21267_ _02998_ _03005_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold571 top_inst.deskew_buff_inst.col_input\[75\] VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[7\] VGND VGND
+ VPWR VPWR net764 sky130_fd_sc_hd__dlygate4sd3_1
X_23006_ top_inst.skew_buff_inst.row\[0\].output_reg\[4\] _04583_ VGND VGND VPWR VPWR
+ _04595_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold593 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[8\] VGND
+ VGND VPWR VPWR net775 sky130_fd_sc_hd__dlygate4sd3_1
X_20218_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _02015_ sky130_fd_sc_hd__buf_2
XFILLER_0_229_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21198_ _02937_ _02938_ _02922_ VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20149_ _01921_ _01957_ _01942_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__a21oi_1
XTAP_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12971_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _05763_ sky130_fd_sc_hd__clkbuf_4
XTAP_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14710_ _07396_ _07397_ _07360_ VGND VGND VPWR VPWR _07399_ sky130_fd_sc_hd__o21ai_1
XTAP_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23908_ clknet_leaf_36_clk _00441_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ net481 _04964_ _04970_ _04968_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__o211a_1
X_15690_ _05311_ VGND VGND VPWR VPWR _08307_ sky130_fd_sc_hd__buf_8
XTAP_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _07329_ _07330_ VGND VGND VPWR VPWR _07331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ net604 _04925_ _04931_ _04929_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23839_ clknet_leaf_89_clk _00372_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_240_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17360_ _09899_ _09900_ VGND VGND VPWR VPWR _09901_ sky130_fd_sc_hd__xnor2_2
X_14572_ _07261_ _07262_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _07264_ sky130_fd_sc_hd__a21o_1
X_11784_ top_inst.axis_out_inst.out_buff_data\[71\] _04890_ VGND VGND VPWR VPWR _04892_
+ sky130_fd_sc_hd__or2_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16311_ _08679_ _08677_ _08686_ _08683_ VGND VGND VPWR VPWR _08893_ sky130_fd_sc_hd__and4_1
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13523_ top_inst.grid_inst.data_path_wires\[2\]\[5\] top_inst.grid_inst.data_path_wires\[2\]\[4\]
+ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__and4_2
X_17291_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[21\] _09631_ VGND
+ VGND VPWR VPWR _09835_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19030_ _11436_ _11437_ _11449_ VGND VGND VPWR VPWR _11451_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16242_ _08824_ _08825_ VGND VGND VPWR VPWR _08826_ sky130_fd_sc_hd__nor2_1
X_13454_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _06212_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12405_ net345 _05243_ _05245_ _05234_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16173_ _08736_ _08738_ VGND VGND VPWR VPWR _08759_ sky130_fd_sc_hd__nand2_1
X_13385_ _06156_ _06157_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15124_ _07771_ _07772_ _07740_ VGND VGND VPWR VPWR _07774_ sky130_fd_sc_hd__a21oi_1
Xoutput109 net109 VGND VGND VPWR VPWR output_tdata[49] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12336_ net678 _05204_ _05206_ _05195_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19932_ _01710_ _01750_ _01752_ _01731_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__a22o_1
X_15055_ _04873_ VGND VGND VPWR VPWR _07707_ sky130_fd_sc_hd__buf_4
XFILLER_0_120_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12267_ net726 _05156_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14006_ _06685_ _06689_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__nor2_1
X_19863_ _01685_ _01686_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__nand2_1
X_12198_ _05127_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__clkbuf_4
Xoutput80 net80 VGND VGND VPWR VPWR output_tdata[22] sky130_fd_sc_hd__clkbuf_4
Xoutput91 net91 VGND VGND VPWR VPWR output_tdata[32] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_207_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18814_ top_inst.grid_inst.data_path_wires\[13\]\[4\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[13\]\[5\]
+ VGND VGND VPWR VPWR _11240_ sky130_fd_sc_hd__a22o_1
XTAP_6070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19794_ _01596_ _01620_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__xor2_1
XTAP_6081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18745_ _11167_ _11172_ _11173_ VGND VGND VPWR VPWR _11175_ sky130_fd_sc_hd__nand3_2
XTAP_5380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15957_ _08565_ _08566_ VGND VGND VPWR VPWR _08567_ sky130_fd_sc_hd__nand2_1
XTAP_5391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14908_ _07558_ _07556_ _07572_ VGND VGND VPWR VPWR _07591_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_163_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18676_ net947 _11116_ net167 VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__o21a_1
XFILLER_0_204_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15888_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[11\] _08374_ VGND
+ VGND VPWR VPWR _08500_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17627_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[5\] _10138_ VGND
+ VGND VPWR VPWR _10139_ sky130_fd_sc_hd__xor2_2
XFILLER_0_118_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14839_ _07450_ _07522_ VGND VGND VPWR VPWR _07524_ sky130_fd_sc_hd__and2_1
XFILLER_0_231_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17558_ _10025_ _10044_ _10042_ _10027_ VGND VGND VPWR VPWR _10073_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16509_ _09040_ _09043_ _09042_ VGND VGND VPWR VPWR _09086_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_188_1358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17489_ top_inst.grid_inst.data_path_wires\[11\]\[0\] VGND VGND VPWR VPWR _10022_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19228_ _11585_ _11615_ _11638_ _11642_ _11637_ VGND VGND VPWR VPWR _11643_ sky130_fd_sc_hd__a32o_1
XFILLER_0_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19159_ _11509_ _11538_ _11536_ VGND VGND VPWR VPWR _11577_ sky130_fd_sc_hd__o21a_1
XFILLER_0_171_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22170_ _03824_ _03829_ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21121_ _02875_ _02869_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21052_ _02814_ _02815_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20003_ _01792_ _01816_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__and2_1
XFILLER_0_236_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21954_ _03630_ _03667_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20905_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[20\] _02559_ _02648_
+ _02675_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_222_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21885_ _03572_ _03583_ _03599_ _03560_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23624_ clknet_leaf_100_clk net511 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_20836_ _02607_ _02609_ VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__xor2_1
XFILLER_0_194_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23555_ clknet_leaf_102_clk _00088_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_20767_ _02542_ _02543_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__and2_1
XFILLER_0_181_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22506_ _04149_ _04160_ _04179_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_190_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23486_ clknet_leaf_138_clk _00019_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[76\]
+ sky130_fd_sc_hd__dfxtp_1
X_20698_ _02463_ _02476_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22437_ _04083_ _04120_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_162_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13170_ _05944_ _05906_ _05947_ _05948_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22368_ _04006_ _04050_ _04051_ _03887_ _04052_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_27_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12121_ net385 _05071_ _05083_ _05075_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__o211a_1
X_24107_ clknet_leaf_14_clk _00640_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_21319_ _03044_ _03056_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22299_ _03950_ _03985_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__xor2_2
XFILLER_0_104_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_236_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24038_ clknet_leaf_42_clk _00571_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_12052_ _04858_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__buf_4
Xhold390 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[9\] VGND
+ VGND VPWR VPWR net572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16860_ _09416_ VGND VGND VPWR VPWR _09417_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1072 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15811_ _08376_ _08379_ VGND VGND VPWR VPWR _08425_ sky130_fd_sc_hd__nor2_1
XFILLER_0_244_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16791_ net170 _09316_ _09348_ _09349_ VGND VGND VPWR VPWR _09350_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18530_ _10990_ _10966_ VGND VGND VPWR VPWR _10992_ sky130_fd_sc_hd__or2b_1
XFILLER_0_232_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15742_ _08355_ _08356_ VGND VGND VPWR VPWR _08357_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_88_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _05750_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11905_ net682 _04951_ _04960_ _04955_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__o211a_1
X_18461_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[10\] _10923_ _10840_
+ VGND VGND VPWR VPWR _10924_ sky130_fd_sc_hd__a21o_1
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15673_ _08287_ _08288_ _08241_ _08243_ VGND VGND VPWR VPWR _08290_ sky130_fd_sc_hd__o211ai_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _05660_ _05670_ _05690_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__a21o_1
XFILLER_0_197_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _09950_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _07313_ VGND VGND VPWR VPWR _07314_ sky130_fd_sc_hd__inv_2
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18392_ _10614_ VGND VGND VPWR VPWR _10857_ sky130_fd_sc_hd__inv_2
X_11836_ net684 _04912_ _04921_ _04916_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _09852_ _09862_ _09883_ _07439_ VGND VGND VPWR VPWR _09885_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14555_ _07205_ _07245_ _07246_ VGND VGND VPWR VPWR _07247_ sky130_fd_sc_hd__nand3_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ top_inst.axis_out_inst.out_buff_data\[64\] _04877_ VGND VGND VPWR VPWR _04882_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_71_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13506_ _06243_ _06256_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__xnor2_1
X_17274_ _09808_ _09810_ _09818_ VGND VGND VPWR VPWR _09819_ sky130_fd_sc_hd__a21o_1
X_14486_ _07178_ _07179_ _07151_ VGND VGND VPWR VPWR _07180_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_99_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_862 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19013_ _11432_ _11433_ VGND VGND VPWR VPWR _11434_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16225_ top_inst.grid_inst.data_path_wires\[8\]\[5\] top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[1\]
+ _08682_ _08676_ VGND VGND VPWR VPWR _08809_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13437_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _06200_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer2 _05265_ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16156_ _08742_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__clkbuf_1
X_13368_ _06140_ _06141_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_224_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15107_ _07621_ top_inst.grid_inst.data_path_wires\[6\]\[5\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[1\]
+ _07626_ VGND VGND VPWR VPWR _07757_ sky130_fd_sc_hd__nand4_1
X_12319_ net941 _05191_ _05197_ _05195_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__o211a_1
X_16087_ _08683_ _08684_ VGND VGND VPWR VPWR _08685_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13299_ _05989_ _06031_ _06074_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_239_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19915_ _01729_ _01730_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__and2b_1
X_15038_ top_inst.grid_inst.data_path_wires\[6\]\[4\] top_inst.grid_inst.data_path_wires\[6\]\[3\]
+ _07629_ _07626_ VGND VGND VPWR VPWR _07690_ sky130_fd_sc_hd__nand4_1
XFILLER_0_227_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19846_ _01642_ _01670_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_235_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16989_ _09505_ _09521_ net214 VGND VGND VPWR VPWR _09543_ sky130_fd_sc_hd__nand3_1
X_19777_ _01488_ _01576_ _01575_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_78_1167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18728_ _11161_ _11150_ VGND VGND VPWR VPWR _11162_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_204_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18659_ _05313_ VGND VGND VPWR VPWR _11116_ sky130_fd_sc_hd__buf_2
XFILLER_0_235_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21670_ _03238_ _03396_ _03397_ _03398_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__o211a_2
XFILLER_0_87_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20621_ _02396_ _02401_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23340_ net161 _04779_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20552_ _02286_ _02293_ _02292_ VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_116_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23271_ net128 _04740_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20483_ _02260_ _02261_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22222_ _03902_ _03910_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__xor2_2
XFILLER_0_15_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22153_ _03842_ _03843_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_242_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21104_ top_inst.grid_inst.data_path_wires\[17\]\[1\] VGND VGND VPWR VPWR _02864_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22084_ net371 _03528_ _03775_ _03776_ _02962_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__o221a_1
XFILLER_0_100_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21035_ _02774_ _02800_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_1212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22986_ net702 _04583_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21937_ _03574_ _03631_ _03651_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__nand3_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _05352_ _05481_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__and2_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21868_ _03584_ _03586_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23607_ clknet_leaf_104_clk net798 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20819_ _02562_ _02588_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__nor2_1
X_24587_ clknet_leaf_20_clk _01120_ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_148_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21799_ _03503_ _03521_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14340_ _05787_ VGND VGND VPWR VPWR _07048_ sky130_fd_sc_hd__buf_4
XFILLER_0_110_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23538_ clknet_leaf_132_clk _00071_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14271_ _06976_ _06981_ VGND VGND VPWR VPWR _06982_ sky130_fd_sc_hd__xnor2_1
X_23469_ clknet_leaf_30_clk _00002_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[123\]
+ sky130_fd_sc_hd__dfxtp_1
X_16010_ _08585_ _08617_ VGND VGND VPWR VPWR _08619_ sky130_fd_sc_hd__and2_1
X_13222_ _05956_ _05958_ _05999_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13153_ _05891_ _05892_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[17\] _05063_
+ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__or2_1
X_13084_ _05750_ top_inst.grid_inst.data_path_wires\[1\]\[5\] _05759_ _05757_ VGND
+ VGND VPWR VPWR _05865_ sky130_fd_sc_hd__and4_1
X_17961_ _10421_ _10423_ _10463_ VGND VGND VPWR VPWR _10465_ sky130_fd_sc_hd__or3_1
XFILLER_0_209_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16912_ _09215_ _09466_ _09467_ VGND VGND VPWR VPWR _09468_ sky130_fd_sc_hd__a21bo_1
X_19700_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[12\] _01480_ VGND
+ VGND VPWR VPWR _01529_ sky130_fd_sc_hd__xnor2_1
X_12035_ _04994_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__buf_2
XFILLER_0_109_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17892_ _10394_ _10396_ VGND VGND VPWR VPWR _10398_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16843_ _09350_ _09398_ _09400_ VGND VGND VPWR VPWR _09401_ sky130_fd_sc_hd__and3_1
X_19631_ _01434_ _01460_ _01461_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__and3_1
XFILLER_0_233_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19562_ _11684_ _11679_ _11709_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__o21a_1
XFILLER_0_233_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16774_ _09207_ _09197_ _09201_ _09203_ VGND VGND VPWR VPWR _09333_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13986_ _06698_ _06699_ VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__or2b_1
XFILLER_0_232_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18513_ _10595_ _10610_ VGND VGND VPWR VPWR _10975_ sky130_fd_sc_hd__nand2_1
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15725_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[7\] _08340_ VGND
+ VGND VPWR VPWR _08341_ sky130_fd_sc_hd__xnor2_1
X_12937_ _04864_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__buf_6
X_19493_ _01279_ _01281_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18444_ _10846_ _10866_ _10864_ VGND VGND VPWR VPWR _10908_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15656_ _08248_ _08254_ VGND VGND VPWR VPWR _08273_ sky130_fd_sc_hd__or2b_1
X_12868_ _05304_ _05641_ _05672_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14607_ _07296_ _07297_ VGND VGND VPWR VPWR _07298_ sky130_fd_sc_hd__xor2_2
XFILLER_0_201_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11819_ _04858_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__buf_4
X_18375_ _10792_ VGND VGND VPWR VPWR _10840_ sky130_fd_sc_hd__clkbuf_4
X_15587_ _08205_ _08206_ VGND VGND VPWR VPWR _08207_ sky130_fd_sc_hd__or2_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _05604_ _05605_ _05538_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__o21a_1
XFILLER_0_185_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17326_ _09853_ _09857_ VGND VGND VPWR VPWR _09868_ sky130_fd_sc_hd__nand2_1
X_14538_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[1\] _07085_ _07089_
+ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _07230_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17257_ _09788_ _09783_ _09801_ VGND VGND VPWR VPWR _09803_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14469_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[1\] _07077_ _07081_
+ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _07163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16208_ _08763_ _08779_ VGND VGND VPWR VPWR _08792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17188_ _09735_ _09736_ VGND VGND VPWR VPWR _09737_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1085 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16139_ _08725_ VGND VGND VPWR VPWR _08726_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_209_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19829_ _01631_ _01640_ _01653_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__a21o_1
XFILLER_0_236_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22840_ top_inst.skew_buff_inst.row\[3\].output_reg\[4\] _03691_ VGND VGND VPWR VPWR
+ _04501_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22771_ _04425_ _04440_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24510_ clknet_leaf_128_clk _01043_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21722_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[19\] _03376_ VGND
+ VGND VPWR VPWR _03448_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_182_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24441_ clknet_leaf_64_clk net904 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[0\].output_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21653_ _03377_ _03381_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20604_ _02344_ _02384_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__or2_1
X_24372_ clknet_leaf_39_clk net407 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].output_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21584_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[13\] _03122_ _03123_
+ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23323_ net153 _04766_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20535_ _02001_ _02015_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[10\]
+ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__and3_1
XFILLER_0_201_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23254_ net120 _04727_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__or2_1
X_20466_ _02248_ _02249_ _02250_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__nand3_2
XFILLER_0_61_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22205_ _03893_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__buf_4
XFILLER_0_28_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23185_ net87 _04687_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20397_ _02181_ _02182_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22136_ _03825_ _03826_ _03688_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[2\]
+ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__and4bb_1
XTAP_6614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22067_ _03758_ _03759_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__nand2_1
XTAP_6669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21018_ _02765_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__inv_2
XTAP_5957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13840_ _06548_ _06551_ _06580_ VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_1075 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_214_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_230_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13771_ _06467_ _06514_ VGND VGND VPWR VPWR _06515_ sky130_fd_sc_hd__xnor2_1
X_22969_ top_inst.skew_buff_inst.row\[1\].output_reg\[4\] _04570_ VGND VGND VPWR VPWR
+ _04574_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15510_ top_inst.grid_inst.data_path_wires\[7\]\[4\] VGND VGND VPWR VPWR _08145_
+ sky130_fd_sc_hd__inv_2
X_12722_ _05530_ _05531_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16490_ _09026_ _09027_ _09067_ VGND VGND VPWR VPWR _09068_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_167_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_214_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15441_ _08076_ _08082_ VGND VGND VPWR VPWR _08083_ sky130_fd_sc_hd__xnor2_1
X_12653_ _05464_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__inv_2
X_24639_ clknet_leaf_25_clk net543 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[115\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_952 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18160_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[2\] _10631_ VGND
+ VGND VPWR VPWR _10632_ sky130_fd_sc_hd__xor2_1
X_15372_ _08013_ _08015_ VGND VGND VPWR VPWR _08016_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12584_ _05372_ _05397_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17111_ _09618_ _09658_ VGND VGND VPWR VPWR _09662_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14323_ _07002_ _07005_ _07031_ VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18091_ _10579_ _04859_ VGND VGND VPWR VPWR _10580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17042_ _09554_ _09556_ net222 VGND VGND VPWR VPWR _09595_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_162_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14254_ _06630_ top_inst.grid_inst.data_path_wires\[3\]\[6\] _06652_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _06965_ sky130_fd_sc_hd__and4b_1
XFILLER_0_0_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13205_ _05933_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__inv_2
X_14185_ top_inst.grid_inst.data_path_wires\[3\]\[7\] _06648_ _06645_ VGND VGND VPWR
+ VPWR _06898_ sky130_fd_sc_hd__and3_2
XFILLER_0_145_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13136_ _05914_ _05915_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ _11343_ _11361_ _11414_ VGND VGND VPWR VPWR _11415_ sky130_fd_sc_hd__a21oi_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13067_ _05840_ _05842_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__or2_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17944_ _10071_ _10445_ _10446_ _10448_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__o211a_1
X_12018_ net795 _05018_ _05025_ _05022_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17875_ _10379_ _10380_ _10038_ _10054_ VGND VGND VPWR VPWR _10381_ sky130_fd_sc_hd__and4b_1
XFILLER_0_40_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19614_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[5\] net195 VGND
+ VGND VPWR VPWR _01445_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16826_ _09375_ _09382_ _09383_ VGND VGND VPWR VPWR _09384_ sky130_fd_sc_hd__nand3_1
XFILLER_0_191_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16757_ _09313_ _09314_ _09315_ VGND VGND VPWR VPWR _09317_ sky130_fd_sc_hd__o21ba_1
X_19545_ _01323_ _01325_ _01376_ _01377_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_177_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13969_ _06686_ _06687_ VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_139_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_139_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_232_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15708_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[6\] _08285_ _08286_
+ VGND VGND VPWR VPWR _08324_ sky130_fd_sc_hd__a21bo_1
X_16688_ _09248_ _09249_ VGND VGND VPWR VPWR _09250_ sky130_fd_sc_hd__nand2_1
X_19476_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[3\]
+ net239 _11696_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__and4_1
XFILLER_0_48_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18427_ _10854_ _10862_ VGND VGND VPWR VPWR _10891_ sky130_fd_sc_hd__or2b_1
X_15639_ _08238_ _08256_ VGND VGND VPWR VPWR _08257_ sky130_fd_sc_hd__xor2_2
XFILLER_0_111_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18358_ _10614_ _10779_ _10823_ VGND VGND VPWR VPWR _10824_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_228_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17309_ _09827_ _09850_ _09851_ VGND VGND VPWR VPWR _09852_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18289_ top_inst.grid_inst.data_path_wires\[12\]\[7\] _10591_ _10600_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _10756_ sky130_fd_sc_hd__nand4_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20320_ _02106_ _02107_ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold901 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[10\] VGND VGND
+ VPWR VPWR net1083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 top_inst.deskew_buff_inst.col_input\[23\] VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[19\] VGND
+ VGND VPWR VPWR net1105 sky130_fd_sc_hd__dlygate4sd3_1
X_20251_ _02040_ _02041_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20182_ _01989_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__buf_4
XFILLER_0_161_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23941_ clknet_leaf_81_clk _00474_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_243_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23872_ clknet_leaf_78_clk _00405_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22823_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[25\] _04488_ _03892_
+ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__a21o_1
XFILLER_0_211_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22754_ _04424_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21705_ _03382_ _03429_ _03411_ _03403_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__a2bb2o_1
X_22685_ _04326_ _04338_ _04357_ _06734_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24424_ clknet_leaf_39_clk net405 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_922 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21636_ _03336_ _03365_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24355_ clknet_leaf_21_clk _00888_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[114\]
+ sky130_fd_sc_hd__dfxtp_1
X_21567_ _03286_ _03298_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__xor2_2
XFILLER_0_244_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_244_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23306_ net145 _04766_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__or2_1
X_20518_ _02299_ _02300_ _02272_ _02273_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21498_ _03197_ _03193_ _03231_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__a21oi_1
X_24286_ clknet_4_4__leaf_clk _00819_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23237_ net112 _04727_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__or2_1
X_20449_ _02232_ net179 VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23168_ _04868_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22119_ _03786_ _03792_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__or2b_1
XFILLER_0_98_1126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23099_ net284 _05323_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__or2_1
X_15990_ _08484_ _08598_ VGND VGND VPWR VPWR _08599_ sky130_fd_sc_hd__xor2_1
XTAP_6455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14941_ _04865_ VGND VGND VPWR VPWR _07611_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17660_ top_inst.grid_inst.data_path_wires\[11\]\[2\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[11\]\[3\]
+ VGND VGND VPWR VPWR _10171_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_215_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14872_ _07548_ VGND VGND VPWR VPWR _07556_ sky130_fd_sc_hd__inv_2
XTAP_5798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16611_ _08870_ _09182_ _09183_ _09184_ VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13823_ _06496_ _06564_ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17591_ _05887_ _10102_ _10103_ _10104_ VGND VGND VPWR VPWR _10105_ sky130_fd_sc_hd__a31o_1
XFILLER_0_214_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16542_ _08679_ _08697_ _08695_ VGND VGND VPWR VPWR _09118_ sky130_fd_sc_hd__and3_1
X_19330_ _11688_ _11677_ VGND VGND VPWR VPWR _11724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13754_ _06492_ _06496_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12705_ _05486_ _05487_ _05515_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__a21oi_4
X_19261_ _05787_ _11674_ _04867_ VGND VGND VPWR VPWR _11675_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_31_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16473_ _09039_ _09015_ _09050_ VGND VGND VPWR VPWR _09051_ sky130_fd_sc_hd__a21o_1
XFILLER_0_168_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13685_ _06385_ _06429_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__and2_1
XFILLER_0_155_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18212_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[4\] _10364_ _10680_
+ _10681_ _09886_ VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__o221a_1
X_15424_ _05353_ VGND VGND VPWR VPWR _08066_ sky130_fd_sc_hd__buf_4
XFILLER_0_156_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12636_ _05447_ _05271_ _05279_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_156_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19192_ _11607_ _11608_ VGND VGND VPWR VPWR _11609_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18143_ _10577_ _10597_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _10617_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15355_ _07956_ _07997_ VGND VGND VPWR VPWR _07999_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12567_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[2\] _05286_ VGND
+ VGND VPWR VPWR _05381_ sky130_fd_sc_hd__and2_1
XFILLER_0_182_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14306_ _06983_ _06982_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__and2b_1
XFILLER_0_123_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18074_ _10536_ _10559_ VGND VGND VPWR VPWR _10574_ sky130_fd_sc_hd__and2b_1
X_15286_ _07886_ _07892_ _07931_ VGND VGND VPWR VPWR _07932_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12498_ _05316_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__clkbuf_16
Xhold208 _00939_ VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17025_ net1040 _09266_ _09577_ _09578_ _07708_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__o221a_1
Xhold219 _00229_ VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ _06905_ _06909_ _06903_ VGND VGND VPWR VPWR _06949_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14168_ _06878_ _06880_ VGND VGND VPWR VPWR _06882_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13119_ _05897_ _05898_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__nand2_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14099_ _06811_ _06813_ VGND VGND VPWR VPWR _06814_ sky130_fd_sc_hd__xnor2_2
X_18976_ _11397_ VGND VGND VPWR VPWR _11398_ sky130_fd_sc_hd__inv_2
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _10377_ _10386_ _10431_ VGND VGND VPWR VPWR _10432_ sky130_fd_sc_hd__a21bo_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_234_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17858_ _06168_ VGND VGND VPWR VPWR _10364_ sky130_fd_sc_hd__buf_4
XFILLER_0_117_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16809_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[7\] _09366_ VGND
+ VGND VPWR VPWR _09367_ sky130_fd_sc_hd__xor2_1
XFILLER_0_178_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17789_ _10295_ _10296_ VGND VGND VPWR VPWR _10297_ sky130_fd_sc_hd__xor2_1
XFILLER_0_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19528_ _01359_ _01360_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19459_ _01291_ _01293_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22470_ _04086_ _04121_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21421_ _03117_ _03156_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24140_ clknet_leaf_144_clk _00673_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_21352_ _02868_ _02893_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20303_ _02088_ _02091_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_188_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24071_ clknet_leaf_84_clk _00604_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_21283_ _02995_ _02996_ _03020_ _03021_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__a211oi_2
Xhold720 top_inst.axis_in_inst.inbuf_bus\[11\] VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold731 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[14\] VGND
+ VGND VPWR VPWR net913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold742 top_inst.deskew_buff_inst.col_input\[73\] VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23022_ _04550_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__buf_4
X_20234_ net737 _01735_ _02026_ _02006_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__o211a_1
Xhold753 top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[1\] VGND VGND
+ VPWR VPWR net935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[17\] VGND VGND
+ VPWR VPWR net946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold775 top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[18\] VGND VGND
+ VPWR VPWR net957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold786 top_inst.deskew_buff_inst.col_input\[17\] VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 top_inst.axis_in_inst.inbuf_bus\[3\] VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20165_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[30\] _01352_ _01524_
+ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20096_ _01884_ _01866_ _01906_ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__and3_1
XTAP_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23924_ clknet_leaf_76_clk _00457_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23855_ clknet_leaf_70_clk _00388_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22806_ _04472_ _04473_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23786_ clknet_leaf_70_clk _00319_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20998_ _02473_ _02743_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22737_ _04377_ _04380_ _04403_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_149_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_1243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13470_ _06186_ _06200_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22668_ _04342_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24407_ clknet_leaf_55_clk net381 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].output_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12421_ net276 _05243_ _05254_ _05247_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21619_ _03322_ _03330_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__nor2_1
XFILLER_0_192_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22599_ _04275_ _04276_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_1126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15140_ _07619_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[2\] _07787_
+ _07788_ VGND VGND VPWR VPWR _07789_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24338_ clknet_leaf_9_clk _00871_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[97\]
+ sky130_fd_sc_hd__dfxtp_1
X_12352_ net306 _05204_ _05215_ _05208_ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15071_ top_inst.grid_inst.data_path_wires\[6\]\[4\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[1\]
+ _07626_ top_inst.grid_inst.data_path_wires\[6\]\[5\] VGND VGND VPWR VPWR _07722_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_1025 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24269_ clknet_leaf_105_clk _00802_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12283_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[30\] _05169_
+ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14022_ _06708_ _06711_ _06712_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__or3_2
XFILLER_0_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18830_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[5\] _09496_ _11254_
+ _11255_ VGND VGND VPWR VPWR _11256_ sky130_fd_sc_hd__a22o_1
XTAP_6230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15973_ _08540_ _08542_ VGND VGND VPWR VPWR _08583_ sky130_fd_sc_hd__or2b_1
X_18761_ _11177_ _11188_ _11189_ _11160_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__o211a_1
XTAP_6285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14924_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[23\] _07595_ VGND
+ VGND VPWR VPWR _07601_ sky130_fd_sc_hd__and2_1
XTAP_5573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17712_ _10220_ _10221_ VGND VGND VPWR VPWR _10222_ sky130_fd_sc_hd__xnor2_1
XTAP_5584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18692_ _10447_ VGND VGND VPWR VPWR _11137_ sky130_fd_sc_hd__buf_2
XFILLER_0_216_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold80 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[20\] VGND
+ VGND VPWR VPWR net262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold91 _00148_ VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14855_ _07538_ _07539_ VGND VGND VPWR VPWR _07540_ sky130_fd_sc_hd__or2_1
XFILLER_0_199_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17643_ _10126_ _10142_ VGND VGND VPWR VPWR _10154_ sky130_fd_sc_hd__nand2_1
XFILLER_0_231_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13806_ _06546_ _06547_ VGND VGND VPWR VPWR _06549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_203_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17574_ top_inst.grid_inst.data_path_wires\[11\]\[1\] top_inst.grid_inst.data_path_wires\[11\]\[0\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _10088_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14786_ _07425_ _07428_ _07471_ _07472_ VGND VGND VPWR VPWR _07473_ sky130_fd_sc_hd__a211o_1
XFILLER_0_202_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11998_ net514 _05010_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16525_ _09053_ _09060_ _09051_ VGND VGND VPWR VPWR _09102_ sky130_fd_sc_hd__o21ai_2
X_19313_ _05269_ _11709_ VGND VGND VPWR VPWR _11710_ sky130_fd_sc_hd__or2_1
X_13737_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[10\] _06242_ _06480_
+ _06481_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_70_clk clknet_4_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16456_ _09000_ _09034_ VGND VGND VPWR VPWR _09035_ sky130_fd_sc_hd__xnor2_1
X_19244_ _11635_ _11658_ VGND VGND VPWR VPWR _11659_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13668_ _06190_ _06212_ VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15407_ _08041_ _08042_ _08048_ VGND VGND VPWR VPWR _08050_ sky130_fd_sc_hd__a21oi_1
X_12619_ _05411_ _05431_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__xnor2_1
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19175_ _11590_ _11591_ VGND VGND VPWR VPWR _11592_ sky130_fd_sc_hd__or2_1
X_16387_ top_inst.grid_inst.data_path_wires\[8\]\[7\] _08693_ _08690_ VGND VGND VPWR
+ VPWR _08967_ sky130_fd_sc_hd__and3_1
XFILLER_0_155_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13599_ _06345_ _06346_ VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18126_ _10604_ _10057_ VGND VGND VPWR VPWR _10605_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15338_ _07950_ _07951_ _07981_ VGND VGND VPWR VPWR _07983_ sky130_fd_sc_hd__or3_1
XFILLER_0_124_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18057_ _10531_ _10532_ _10557_ VGND VGND VPWR VPWR _10558_ sky130_fd_sc_hd__a21oi_1
X_15269_ _07913_ _07914_ VGND VGND VPWR VPWR _07915_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17008_ _09553_ _09560_ _09561_ VGND VGND VPWR VPWR _09562_ sky130_fd_sc_hd__or3_4
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_223_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18959_ _11381_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21970_ top_inst.grid_inst.data_path_wires\[18\]\[1\] VGND VGND VPWR VPWR _03682_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_207_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer12 net193 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_1
Xrebuffer23 _07059_ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_1
XFILLER_0_179_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20921_ _02688_ _02689_ _02466_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__a21oi_1
Xrebuffer34 _09205_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_221_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer45 _09205_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer56 _01462_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer67 _01401_ VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23640_ clknet_leaf_126_clk net403 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20852_ _02528_ _02616_ _02623_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__nand3_1
Xrebuffer78 _07151_ VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_166_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_230_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23571_ clknet_leaf_107_clk _00104_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20783_ _02468_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_61_clk clknet_4_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22522_ _04193_ _04202_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__xor2_1
XFILLER_0_190_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22453_ _04135_ _03695_ _04104_ _04100_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_49_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21404_ _03138_ _03139_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22384_ _03711_ top_inst.grid_inst.data_path_wires\[18\]\[6\] VGND VGND VPWR VPWR
+ _04069_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24123_ clknet_leaf_11_clk _00656_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_32_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21335_ _03064_ _03065_ _03071_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__a21o_2
XFILLER_0_241_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24054_ clknet_leaf_34_clk _00587_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_241_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold550 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[0\]\[0\] VGND VGND
+ VPWR VPWR net732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21266_ _02999_ _03004_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__xor2_1
Xhold561 top_inst.axis_out_inst.out_buff_data\[74\] VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold572 _00050_ VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 _00933_ VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__dlygate4sd3_1
X_23005_ net979 _04588_ _04594_ _04590_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20217_ _01995_ _11163_ _02014_ _02006_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold594 top_inst.axis_out_inst.out_buff_data\[64\] VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__dlygate4sd3_1
X_21197_ _02922_ _02937_ _02938_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__or3_1
XFILLER_0_204_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20148_ _01950_ _01958_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_244_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_205_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20079_ _01562_ _01892_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__nor2_1
X_12970_ _05741_ _05756_ _05762_ _05743_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__o211a_1
XTAP_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23907_ clknet_leaf_37_clk _00440_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ top_inst.axis_out_inst.out_buff_data\[34\] _04969_ VGND VGND VPWR VPWR _04970_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_197_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _07079_ _07074_ _07082_ _07086_ VGND VGND VPWR VPWR _07330_ sky130_fd_sc_hd__nand4_1
XTAP_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ net348 _04930_ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__or2_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23838_ clknet_leaf_89_clk _00371_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[7\] _07261_ _07262_
+ VGND VGND VPWR VPWR _07263_ sky130_fd_sc_hd__nand3_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23769_ clknet_leaf_66_clk _00302_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11783_ net360 _04885_ _04891_ _04889_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__o211a_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_52_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16310_ _08889_ _08891_ VGND VGND VPWR VPWR _08892_ sky130_fd_sc_hd__xnor2_1
X_13522_ top_inst.grid_inst.data_path_wires\[2\]\[2\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[2\]
+ _06253_ _06252_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[4\] VGND
+ VGND VPWR VPWR _06272_ sky130_fd_sc_hd__a32o_1
X_17290_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[20\] _09628_ _09629_
+ VGND VGND VPWR VPWR _09834_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16241_ _08822_ _08823_ _08791_ VGND VGND VPWR VPWR _08825_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13453_ _06190_ _06204_ _06211_ _06207_ VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12404_ net341 _05235_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__or2_1
X_16172_ _08755_ _08757_ VGND VGND VPWR VPWR _08758_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13384_ _06155_ _06146_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15123_ _07740_ _07771_ _07772_ VGND VGND VPWR VPWR _07773_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12335_ net292 _05196_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_1183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19931_ _01718_ _01716_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__nand2_1
X_15054_ _07703_ _07704_ _07057_ VGND VGND VPWR VPWR _07706_ sky130_fd_sc_hd__a21o_1
XFILLER_0_220_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12266_ net825 _05164_ _05166_ _05155_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14005_ _06707_ _06722_ VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__xor2_1
XFILLER_0_107_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19862_ _01683_ _01684_ _01527_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput70 net70 VGND VGND VPWR VPWR output_tdata[13] sky130_fd_sc_hd__clkbuf_4
X_12197_ _04873_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__buf_2
Xoutput81 net81 VGND VGND VPWR VPWR output_tdata[23] sky130_fd_sc_hd__clkbuf_4
X_18813_ _11217_ _11220_ _11218_ VGND VGND VPWR VPWR _11239_ sky130_fd_sc_hd__o21ai_2
Xoutput92 net92 VGND VGND VPWR VPWR output_tdata[33] sky130_fd_sc_hd__clkbuf_4
XTAP_6060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19793_ _01597_ _01619_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__xnor2_1
XTAP_6082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18744_ _11172_ _11173_ _11167_ VGND VGND VPWR VPWR _11174_ sky130_fd_sc_hd__a21o_1
XFILLER_0_207_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15956_ _08484_ _08564_ VGND VGND VPWR VPWR _08566_ sky130_fd_sc_hd__or2_1
XTAP_5381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14907_ _07570_ _07589_ VGND VGND VPWR VPWR _07590_ sky130_fd_sc_hd__xnor2_1
X_18675_ net939 _11116_ net167 VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__o21a_1
X_15887_ _08152_ _08159_ _08445_ _08444_ _08150_ VGND VGND VPWR VPWR _08499_ sky130_fd_sc_hd__a32o_1
XTAP_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17626_ _10136_ _10137_ VGND VGND VPWR VPWR _10138_ sky130_fd_sc_hd__nand2_1
X_14838_ _07450_ _07522_ VGND VGND VPWR VPWR _07523_ sky130_fd_sc_hd__nor2_1
XFILLER_0_188_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14769_ _07421_ _07422_ VGND VGND VPWR VPWR _07456_ sky130_fd_sc_hd__or2b_1
XFILLER_0_188_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17557_ _10022_ _10047_ VGND VGND VPWR VPWR _10072_ sky130_fd_sc_hd__nand2_1
XFILLER_0_175_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16508_ _09040_ _09084_ VGND VGND VPWR VPWR _09085_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17488_ net989 _08183_ _10021_ _09231_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19227_ _11620_ _11618_ VGND VGND VPWR VPWR _11642_ sky130_fd_sc_hd__nand2_1
X_16439_ _09003_ _09004_ _09017_ VGND VGND VPWR VPWR _09018_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19158_ _11550_ _11575_ VGND VGND VPWR VPWR _11576_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18109_ _10592_ _08674_ VGND VGND VPWR VPWR _10593_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19089_ _11470_ _11475_ _11473_ VGND VGND VPWR VPWR _11508_ sky130_fd_sc_hd__a21o_1
XFILLER_0_164_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21120_ top_inst.grid_inst.data_path_wires\[17\]\[6\] VGND VGND VPWR VPWR _02875_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21051_ _02814_ _02815_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20002_ _07057_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__buf_4
XFILLER_0_226_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_213_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21953_ _03628_ _03666_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_193_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20904_ _02674_ _02647_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21884_ _03601_ _03602_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_234_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23623_ clknet_leaf_100_clk net470 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20835_ _02581_ _02608_ VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__nand2_1
XFILLER_0_178_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_34_clk clknet_4_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23554_ clknet_leaf_129_clk _00087_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20766_ _02535_ _02541_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__nand2_1
XFILLER_0_175_871 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22505_ _04154_ _04184_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23485_ clknet_leaf_138_clk _00018_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[75\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20697_ _02464_ _02475_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__xor2_1
XFILLER_0_220_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22436_ _04118_ _04119_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22367_ _04013_ _04012_ _04045_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_32_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24106_ clknet_leaf_115_clk _00639_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_2
X_12120_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[24\] _05076_
+ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21318_ _03049_ _03055_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__xor2_1
XFILLER_0_237_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22298_ _03693_ _03983_ _03984_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_102_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24037_ clknet_leaf_42_clk _00570_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_12051_ net477 _05031_ _05043_ _05035_ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold380 _00068_ VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__dlygate4sd3_1
X_21249_ _02963_ _02987_ _10831_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__o21a_1
XFILLER_0_229_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold391 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[16\] VGND
+ VGND VPWR VPWR net573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_1084 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15810_ _08421_ _08423_ VGND VGND VPWR VPWR _08424_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_244_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16790_ _09346_ _09347_ _09300_ _09302_ VGND VGND VPWR VPWR _09349_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_102_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_244_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15741_ _08143_ _08167_ VGND VGND VPWR VPWR _08356_ sky130_fd_sc_hd__nand2_2
X_12953_ top_inst.grid_inst.data_path_wires\[1\]\[6\] VGND VGND VPWR VPWR _05750_
+ sky130_fd_sc_hd__buf_2
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11904_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[27\] _04956_
+ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__or2_1
X_18460_ _10793_ VGND VGND VPWR VPWR _10923_ sky130_fd_sc_hd__clkbuf_4
X_15672_ _08241_ _08243_ _08287_ _08288_ VGND VGND VPWR VPWR _08289_ sky130_fd_sc_hd__a211o_1
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12884_ _05655_ _05689_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14623_ _07272_ _07305_ VGND VGND VPWR VPWR _07313_ sky130_fd_sc_hd__nand2_1
X_17411_ _09661_ _09949_ VGND VGND VPWR VPWR _09950_ sky130_fd_sc_hd__and2_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18391_ top_inst.grid_inst.data_path_wires\[12\]\[2\] _10614_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[6\]
+ top_inst.grid_inst.data_path_wires\[12\]\[3\] VGND VGND VPWR VPWR _10856_ sky130_fd_sc_hd__and4b_1
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11835_ top_inst.axis_out_inst.out_buff_data\[93\] _04917_ VGND VGND VPWR VPWR _04921_
+ sky130_fd_sc_hd__or2_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clknet_4_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17342_ _09852_ _09862_ _09883_ VGND VGND VPWR VPWR _09884_ sky130_fd_sc_hd__a21oi_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[5\] _07069_ _07243_
+ _07244_ VGND VGND VPWR VPWR _07246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_200_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ net499 _04860_ _04881_ _04875_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13505_ _06250_ _06255_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__xor2_1
X_17273_ _09812_ _09817_ VGND VGND VPWR VPWR _09818_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14485_ _07169_ _07170_ _07177_ VGND VGND VPWR VPWR _07179_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16224_ _08767_ _08768_ _08766_ VGND VGND VPWR VPWR _08808_ sky130_fd_sc_hd__o21a_1
X_19012_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[10\] _11340_ VGND
+ VGND VPWR VPWR _11433_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13436_ _05753_ _06192_ _06199_ _06183_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer3 _05265_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16155_ _08197_ _08741_ VGND VGND VPWR VPWR _08742_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13367_ _06106_ _06109_ _06138_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15106_ top_inst.grid_inst.data_path_wires\[6\]\[5\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[1\]
+ _07626_ top_inst.grid_inst.data_path_wires\[6\]\[6\] VGND VGND VPWR VPWR _07756_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12318_ net449 _05196_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16086_ _05772_ VGND VGND VPWR VPWR _08684_ sky130_fd_sc_hd__buf_2
X_13298_ _06028_ _06030_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15037_ top_inst.grid_inst.data_path_wires\[6\]\[3\] top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[1\]
+ _07626_ top_inst.grid_inst.data_path_wires\[6\]\[4\] VGND VGND VPWR VPWR _07689_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19914_ _05787_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__buf_4
X_12249_ net483 _05151_ _05157_ _05155_ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19845_ _01654_ _01669_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19776_ _01600_ _01602_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__xor2_1
XFILLER_0_208_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16988_ _09501_ _09504_ _09541_ VGND VGND VPWR VPWR _09542_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_235_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18727_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[5\] VGND VGND
+ VPWR VPWR _11161_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_190_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15939_ _08477_ _08511_ VGND VGND VPWR VPWR _08550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18658_ _10071_ _11114_ _11115_ _10620_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__o211a_1
XFILLER_0_231_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_235_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_203_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17609_ _10099_ _10102_ VGND VGND VPWR VPWR _10122_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18589_ _11044_ _11048_ VGND VGND VPWR VPWR _11049_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_clk clknet_4_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20620_ _02399_ _02400_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20551_ _02327_ _02333_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23270_ net622 _04739_ _04747_ _04743_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__o211a_1
X_20482_ net871 _01735_ _02266_ _02035_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22221_ _03907_ _03909_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__xor2_2
XFILLER_0_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_242_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22152_ _03751_ _03773_ _03798_ _03802_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__o31a_1
XFILLER_0_219_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21103_ _01987_ _11142_ _02863_ _02707_ VGND VGND VPWR VPWR _00806_ sky130_fd_sc_hd__o211a_1
XFILLER_0_242_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22083_ _03773_ _03774_ _07595_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21034_ _02798_ _02799_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_227_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_1072 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22985_ _04863_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_215_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21936_ _03574_ _03631_ _03651_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21867_ _03584_ _03586_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__nor2_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23606_ clknet_leaf_104_clk _00139_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20818_ _02568_ _02592_ _04870_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__o21a_1
X_24586_ clknet_leaf_141_clk _01119_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_132_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21798_ _03519_ _03520_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__and2_1
XFILLER_0_231_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23537_ clknet_leaf_141_clk _00070_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20749_ _02518_ _02525_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_231_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14270_ _06980_ VGND VGND VPWR VPWR _06981_ sky130_fd_sc_hd__inv_2
X_23468_ clknet_leaf_30_clk _00001_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[122\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13221_ _05953_ _05955_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22419_ _04067_ _04102_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23399_ net63 _04658_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13152_ _05929_ _05930_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12103_ net573 _05071_ _05073_ _05062_ VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__o211a_1
XFILLER_0_237_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13083_ _05824_ _05827_ _05825_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__a21bo_1
X_17960_ _10421_ _10423_ _10463_ VGND VGND VPWR VPWR _10464_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218_842 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16911_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[4\] _09209_ net203
+ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _09467_ sky130_fd_sc_hd__a22o_1
X_12034_ net1105 _05023_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__or2_1
X_17891_ _10394_ _10396_ VGND VGND VPWR VPWR _10397_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19630_ net196 _01459_ _01418_ _01435_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_205_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16842_ _09399_ _09397_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _09400_ sky130_fd_sc_hd__a21o_1
XFILLER_0_217_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19561_ _01357_ _01374_ _01375_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__nand3_1
XFILLER_0_205_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_189_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16773_ _09329_ _09330_ _09324_ VGND VGND VPWR VPWR _09332_ sky130_fd_sc_hd__a21o_1
X_13985_ _06703_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18512_ _10967_ _10973_ VGND VGND VPWR VPWR _10974_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_232_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12936_ top_inst.grid_inst.data_path_wires\[1\]\[1\] VGND VGND VPWR VPWR _05738_
+ sky130_fd_sc_hd__clkbuf_4
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15724_ _08338_ _08339_ VGND VGND VPWR VPWR _08340_ sky130_fd_sc_hd__xnor2_1
X_19492_ _01323_ _01324_ _01306_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__a21o_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18443_ _10889_ _10906_ VGND VGND VPWR VPWR _10907_ sky130_fd_sc_hd__xnor2_1
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12867_ _05304_ _05641_ _05672_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__a21oi_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15655_ _08253_ _08249_ VGND VGND VPWR VPWR _08272_ sky130_fd_sc_hd__or2b_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14606_ _07243_ _07245_ VGND VGND VPWR VPWR _07297_ sky130_fd_sc_hd__and2_1
XFILLER_0_205_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11818_ net474 _04898_ _04910_ _04902_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18374_ _10837_ _10838_ VGND VGND VPWR VPWR _10839_ sky130_fd_sc_hd__nand2_1
X_15586_ _08203_ _08204_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[3\]
+ VGND VGND VPWR VPWR _08206_ sky130_fd_sc_hd__a21oi_1
X_12798_ _05538_ _05604_ _05605_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__nor3_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[0\] _07085_ _07089_
+ VGND VGND VPWR VPWR _07229_ sky130_fd_sc_hd__and3_1
X_17325_ _09858_ _09859_ VGND VGND VPWR VPWR _09867_ sky130_fd_sc_hd__or2b_1
XFILLER_0_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11749_ net777 _04860_ _04866_ _04870_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14468_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[4\] _07136_ _07137_
+ VGND VGND VPWR VPWR _07162_ sky130_fd_sc_hd__a21bo_1
X_17256_ _09788_ _09783_ _09801_ VGND VGND VPWR VPWR _09802_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16207_ _08784_ _08783_ VGND VGND VPWR VPWR _08791_ sky130_fd_sc_hd__nor2_1
X_13419_ _05741_ _05256_ _06187_ _06183_ VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__o211a_1
X_17187_ _09678_ _09733_ _09734_ VGND VGND VPWR VPWR _09736_ sky130_fd_sc_hd__and3_1
X_14399_ _07066_ _07062_ _07061_ _07065_ VGND VGND VPWR VPWR _07097_ sky130_fd_sc_hd__nand4_1
XFILLER_0_10_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16138_ _08690_ _08688_ _08664_ _08661_ VGND VGND VPWR VPWR _08725_ sky130_fd_sc_hd__and4_2
XFILLER_0_45_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16069_ top_inst.grid_inst.data_path_wires\[8\]\[4\] VGND VGND VPWR VPWR _08671_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_clk clknet_4_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19828_ _01637_ _01639_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__and2_1
XFILLER_0_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_235_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19759_ _01585_ _01586_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__nor2_2
XFILLER_0_196_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22770_ _04438_ _04439_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_231_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21721_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[18\] _03421_ _03422_
+ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_8_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_231_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24440_ clknet_leaf_54_clk _00973_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21652_ _03379_ _03380_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20603_ _02343_ _02381_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_975 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24371_ clknet_leaf_37_clk net656 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].output_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21583_ _03279_ _03282_ _03284_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_7_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23322_ net657 _04765_ _04776_ _04769_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20534_ _02001_ _02015_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[10\]
+ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_160_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23253_ net1025 _04726_ _04737_ _04730_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20465_ _02191_ _02198_ _02197_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_63_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22204_ _03891_ _03892_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23184_ net749 _04685_ _04698_ _04691_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20396_ _01986_ _02178_ _02179_ _02180_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__nor4_1
XFILLER_0_113_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22135_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[3\]
+ top_inst.grid_inst.data_path_wires\[18\]\[3\] top_inst.grid_inst.data_path_wires\[18\]\[2\]
+ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__and4_1
XTAP_6604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22066_ _03688_ _03686_ _03700_ _03697_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__nand4_1
XTAP_6659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21017_ _02778_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__inv_2
XFILLER_0_215_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_214_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_214_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_230_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13770_ _06512_ _06513_ VGND VGND VPWR VPWR _06514_ sky130_fd_sc_hd__nor2_1
X_22968_ net702 _04562_ _04573_ _04564_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12721_ _05298_ _05292_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21919_ _03634_ _03628_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__or2b_1
XFILLER_0_74_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22899_ net394 _04530_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15440_ _08077_ _08081_ VGND VGND VPWR VPWR _08082_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_214_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12652_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[0\]
+ _05300_ _05305_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__and4_1
XFILLER_0_194_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24638_ clknet_leaf_21_clk _01171_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[114\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15371_ _07971_ _07974_ _08014_ VGND VGND VPWR VPWR _08015_ sky130_fd_sc_hd__a21bo_1
X_12583_ _05394_ _05396_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__xnor2_1
X_24569_ clknet_leaf_141_clk _01102_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_136_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_1112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14322_ _06936_ _07030_ VGND VGND VPWR VPWR _07031_ sky130_fd_sc_hd__xnor2_1
X_17110_ _04873_ VGND VGND VPWR VPWR _09661_ sky130_fd_sc_hd__buf_4
XFILLER_0_110_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18090_ top_inst.grid_inst.data_path_wires\[12\]\[1\] VGND VGND VPWR VPWR _10579_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_167_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17041_ _09590_ _09593_ VGND VGND VPWR VPWR _09594_ sky130_fd_sc_hd__xor2_1
XFILLER_0_163_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14253_ _06652_ top_inst.grid_inst.data_path_wires\[3\]\[6\] _06630_ _06963_ VGND
+ VGND VPWR VPWR _06964_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_80_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1056 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13204_ _05976_ _05981_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__xor2_1
X_14184_ _06895_ _06896_ VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13135_ _05832_ _05870_ _05868_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__a21o_1
XFILLER_0_238_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18992_ _11360_ _11358_ VGND VGND VPWR VPWR _11414_ sky130_fd_sc_hd__and2b_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1054 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13066_ _05847_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__clkbuf_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _10447_ VGND VGND VPWR VPWR _10448_ sky130_fd_sc_hd__buf_4
XFILLER_0_225_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12017_ net563 _05023_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__or2_1
X_17874_ _10378_ _10059_ _10056_ top_inst.grid_inst.data_path_wires\[11\]\[5\] VGND
+ VGND VPWR VPWR _10380_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_1252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19613_ _01402_ _01443_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__xor2_1
XFILLER_0_217_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16825_ _09380_ _09381_ _09338_ VGND VGND VPWR VPWR _09383_ sky130_fd_sc_hd__a21o_1
XFILLER_0_233_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_232_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19544_ _01374_ _01375_ _01357_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_233_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16756_ net170 _09314_ _09315_ VGND VGND VPWR VPWR _09316_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_152_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13968_ top_inst.grid_inst.data_path_wires\[3\]\[3\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[3\]\[4\]
+ VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15707_ _08310_ _08322_ VGND VGND VPWR VPWR _08323_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_232_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12919_ _05703_ _05701_ _05608_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19475_ _11697_ _11692_ _11696_ _11693_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__a22oi_1
X_16687_ _09194_ _09188_ _09197_ _09202_ VGND VGND VPWR VPWR _09249_ sky130_fd_sc_hd__nand4_1
X_13899_ top_inst.grid_inst.data_path_wires\[3\]\[6\] VGND VGND VPWR VPWR _06632_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_236_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18426_ _10861_ _10860_ VGND VGND VPWR VPWR _10890_ sky130_fd_sc_hd__or2b_1
XFILLER_0_174_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15638_ _08247_ _08255_ VGND VGND VPWR VPWR _08256_ sky130_fd_sc_hd__xor2_2
XFILLER_0_111_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18357_ _10778_ _10777_ VGND VGND VPWR VPWR _10823_ sky130_fd_sc_hd__and2b_1
XFILLER_0_145_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15569_ _08135_ _08159_ VGND VGND VPWR VPWR _08190_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17308_ _09819_ _09830_ _09846_ VGND VGND VPWR VPWR _09851_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18288_ _10591_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[0\]
+ top_inst.grid_inst.data_path_wires\[12\]\[7\] VGND VGND VPWR VPWR _10755_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17239_ _09661_ _09785_ VGND VGND VPWR VPWR _09786_ sky130_fd_sc_hd__and2_1
XFILLER_0_181_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold902 top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[9\] VGND VGND
+ VPWR VPWR net1084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 top_inst.deskew_buff_inst.col_input\[21\] VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20250_ _02037_ _02038_ _02039_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__and3_1
Xhold924 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[12\] VGND
+ VGND VPWR VPWR net1106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20181_ top_inst.grid_inst.data_path_wires\[16\]\[1\] VGND VGND VPWR VPWR _01989_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23940_ clknet_leaf_81_clk _00473_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23871_ clknet_leaf_78_clk _00404_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22822_ _03700_ _03698_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22753_ _07707_ _04423_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21704_ _03420_ _03430_ VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__xor2_1
XFILLER_0_176_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22684_ _04326_ _04338_ _04357_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_165_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24423_ clknet_leaf_56_clk _00956_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21635_ _03362_ _03364_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__xor2_2
XFILLER_0_192_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24354_ clknet_leaf_26_clk _00887_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[113\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21566_ _03295_ _03297_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_244_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23305_ net927 _04765_ _04767_ _04756_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__o211a_1
XFILLER_0_244_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20517_ _02272_ _02273_ _02299_ _02300_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_105_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24285_ clknet_leaf_10_clk _00818_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_244_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21497_ _03198_ _03230_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23236_ net796 _04726_ _04728_ _04717_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20448_ _01990_ _02229_ _02230_ _02231_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__nor4_1
XFILLER_0_244_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23167_ net79 _04687_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__or2_1
XTAP_6401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20379_ _02164_ _02165_ _02104_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_101_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22118_ _03791_ _03787_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__or2b_1
XFILLER_0_98_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23098_ net624 _10541_ _04647_ _04643_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__o211a_1
XTAP_6456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_238_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14940_ top_inst.grid_inst.data_path_wires\[6\]\[2\] VGND VGND VPWR VPWR _07610_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22049_ _03684_ _03700_ _03698_ _03686_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__a22o_1
XFILLER_0_237_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14871_ net1062 _06660_ _07555_ _07092_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16610_ _07617_ VGND VGND VPWR VPWR _09184_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_187_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13822_ _06562_ _06563_ VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__and2_1
X_17590_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[3\] _05730_ VGND
+ VGND VPWR VPWR _10104_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16541_ _09086_ _09085_ VGND VGND VPWR VPWR _09117_ sky130_fd_sc_hd__or2b_1
X_13753_ _06492_ _06496_ VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12704_ _05505_ _05514_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__xnor2_2
X_19260_ _11643_ _11659_ _11672_ _11673_ VGND VGND VPWR VPWR _11674_ sky130_fd_sc_hd__a211o_1
X_16472_ _09048_ _09049_ VGND VGND VPWR VPWR _09050_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13684_ _06385_ _06429_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18211_ _10678_ _10679_ _09292_ VGND VGND VPWR VPWR _10681_ sky130_fd_sc_hd__a21o_1
X_12635_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _05447_ sky130_fd_sc_hd__inv_2
XFILLER_0_182_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15423_ _08029_ _08065_ _05440_ VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19191_ _11606_ _11588_ VGND VGND VPWR VPWR _11608_ sky130_fd_sc_hd__or2b_1
XFILLER_0_2_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15354_ _07956_ _07997_ VGND VGND VPWR VPWR _07998_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18142_ _05787_ VGND VGND VPWR VPWR _10616_ sky130_fd_sc_hd__buf_4
XFILLER_0_109_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12566_ _05378_ _05379_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14305_ _06995_ _07014_ VGND VGND VPWR VPWR _07015_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15285_ _07885_ _07883_ VGND VGND VPWR VPWR _07931_ sky130_fd_sc_hd__and2b_1
X_18073_ _10564_ _10572_ VGND VGND VPWR VPWR _10573_ sky130_fd_sc_hd__xnor2_1
X_12497_ _05315_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__buf_6
XFILLER_0_0_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14236_ _06943_ _06947_ VGND VGND VPWR VPWR _06948_ sky130_fd_sc_hd__xnor2_1
X_17024_ _09540_ _09535_ _09576_ _07439_ VGND VGND VPWR VPWR _09578_ sky130_fd_sc_hd__a31o_1
Xhold209 top_inst.axis_out_inst.out_buff_data\[85\] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_238_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1020 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14167_ _06878_ _06880_ VGND VGND VPWR VPWR _06881_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _05748_ _05761_ _05895_ _05896_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__nand4_2
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _06770_ _06771_ _06812_ VGND VGND VPWR VPWR _06813_ sky130_fd_sc_hd__o21ba_1
X_18975_ top_inst.grid_inst.data_path_wires\[13\]\[6\] top_inst.grid_inst.data_path_wires\[13\]\[5\]
+ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _11397_ sky130_fd_sc_hd__and4_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13049_ top_inst.grid_inst.data_path_wires\[1\]\[2\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[2\]
+ _05812_ _05811_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[4\] VGND
+ VGND VPWR VPWR _05831_ sky130_fd_sc_hd__a32o_1
X_17926_ _10381_ _10383_ _10385_ VGND VGND VPWR VPWR _10431_ sky130_fd_sc_hd__or3_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17857_ _10071_ _10362_ _10363_ _10049_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__o211a_1
XFILLER_0_234_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16808_ _09364_ _09365_ VGND VGND VPWR VPWR _09366_ sky130_fd_sc_hd__nand2_1
X_17788_ _10040_ _10047_ VGND VGND VPWR VPWR _10296_ sky130_fd_sc_hd__nand2_4
XFILLER_0_89_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19527_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[3\]
+ _11695_ net195 VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__and4_1
X_16739_ _09296_ _09297_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[5\]
+ VGND VGND VPWR VPWR _09299_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19458_ _01250_ _01251_ _01292_ _01256_ VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18409_ _10871_ _10873_ VGND VGND VPWR VPWR _10874_ sky130_fd_sc_hd__nor2_1
X_19389_ _01223_ _01224_ _09292_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21420_ _03154_ _03155_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21351_ _03086_ _03087_ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20302_ _02089_ _02090_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__or2_2
X_24070_ clknet_leaf_84_clk _00603_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_114_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold710 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[5\] VGND
+ VGND VPWR VPWR net892 sky130_fd_sc_hd__dlygate4sd3_1
X_21282_ _03018_ _03019_ _02997_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__a21oi_1
Xhold721 top_inst.axis_in_inst.inbuf_bus\[0\] VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold732 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[20\] VGND
+ VGND VPWR VPWR net914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23021_ net983 _04603_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__or2_1
XFILLER_0_163_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20233_ _02024_ _02025_ _08181_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__o21ai_1
Xhold743 top_inst.deskew_buff_inst.col_input\[20\] VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[2\]\[0\] VGND VGND
+ VPWR VPWR net936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold765 top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[20\] VGND VGND
+ VPWR VPWR net947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 top_inst.deskew_buff_inst.col_input\[21\] VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold787 top_inst.axis_in_inst.inbuf_bus\[10\] VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold798 _00977_ VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__dlygate4sd3_1
X_20164_ _01961_ _01973_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20095_ net1098 _01202_ _01907_ _01908_ _01863_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__o221a_1
XTAP_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23923_ clknet_leaf_76_clk _00456_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23854_ clknet_leaf_69_clk _00387_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22805_ _04471_ _04467_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__or2b_1
XFILLER_0_135_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23785_ clknet_leaf_65_clk _00318_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20997_ _02751_ _02752_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__nand2_1
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22736_ _04382_ _04404_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22667_ _07707_ _04341_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24406_ clknet_leaf_57_clk net390 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].output_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12420_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[25\] _05248_
+ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__or2_1
X_21618_ _03315_ _03319_ _03317_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22598_ _04273_ _04274_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__and2_1
XFILLER_0_168_1176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_7__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_4_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24337_ clknet_leaf_9_clk _00870_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[96\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12351_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[27\] _05209_
+ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21549_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[12\] _03122_ _03123_
+ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15070_ _07610_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.weight_reg\[2\] _07697_
+ _07670_ _07635_ VGND VGND VPWR VPWR _07721_ sky130_fd_sc_hd__a32o_1
XFILLER_0_161_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24268_ clknet_leaf_100_clk _00801_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_12282_ net790 _05164_ _05175_ _05168_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_1195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14021_ _06737_ _06721_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__nor2_1
X_23219_ net103 _04714_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24199_ clknet_leaf_116_clk _00732_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_6220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18760_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[2\] _10639_ VGND
+ VGND VPWR VPWR _11189_ sky130_fd_sc_hd__or2_1
XTAP_6275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15972_ _08580_ _08581_ VGND VGND VPWR VPWR _08582_ sky130_fd_sc_hd__xnor2_1
XTAP_6286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17711_ _10180_ _10182_ VGND VGND VPWR VPWR _10221_ sky130_fd_sc_hd__nor2_1
X_14923_ _07593_ _07600_ _07594_ VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__o21a_1
XTAP_5563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18691_ _11135_ _11133_ VGND VGND VPWR VPWR _11136_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold81 _00155_ VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold92 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[26\] VGND
+ VGND VPWR VPWR net274 sky130_fd_sc_hd__dlygate4sd3_1
X_17642_ _10153_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__clkbuf_1
X_14854_ _07492_ _07507_ _07505_ VGND VGND VPWR VPWR _07539_ sky130_fd_sc_hd__o21a_1
XFILLER_0_188_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13805_ _06546_ _06547_ VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__or2_1
X_17573_ _10022_ _10050_ _10047_ _10025_ VGND VGND VPWR VPWR _10087_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14785_ _07455_ _07469_ VGND VGND VPWR VPWR _07472_ sky130_fd_sc_hd__and2_1
X_11997_ net779 _05004_ _05013_ _05008_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_230_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19312_ _11708_ VGND VGND VPWR VPWR _11709_ sky130_fd_sc_hd__clkbuf_4
X_16524_ _09099_ _09100_ VGND VGND VPWR VPWR _09101_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13736_ _06447_ _06443_ _06479_ _06404_ VGND VGND VPWR VPWR _06481_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_97_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19243_ _11655_ _11657_ VGND VGND VPWR VPWR _11658_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16455_ _09032_ _09033_ VGND VGND VPWR VPWR _09034_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13667_ _06411_ _06412_ VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15406_ _08041_ _08042_ _08048_ VGND VGND VPWR VPWR _08049_ sky130_fd_sc_hd__and3_1
X_12618_ _05422_ _05430_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__xnor2_1
X_19174_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[14\] _11469_ VGND
+ VGND VPWR VPWR _11591_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16386_ _08964_ _08965_ VGND VGND VPWR VPWR _08966_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13598_ _06342_ _06344_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18125_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _10604_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12549_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[4\] _05271_ _05278_
+ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _05364_ sky130_fd_sc_hd__a22o_1
X_15337_ _07950_ _07951_ _07981_ VGND VGND VPWR VPWR _07982_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_26_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18056_ _10533_ _10522_ VGND VGND VPWR VPWR _10557_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1 _02869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15268_ _07871_ _07873_ _07870_ VGND VGND VPWR VPWR _07914_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17007_ _09557_ _09558_ net1121 VGND VGND VPWR VPWR _09561_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_160_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14219_ _06891_ _06894_ _06892_ VGND VGND VPWR VPWR _06931_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_112_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15199_ _07788_ _07790_ _07846_ VGND VGND VPWR VPWR _07847_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_238_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18958_ _10641_ _11380_ VGND VGND VPWR VPWR _11381_ sky130_fd_sc_hd__and2_1
XFILLER_0_225_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17909_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[12\] _10236_ VGND
+ VGND VPWR VPWR _10414_ sky130_fd_sc_hd__xnor2_1
X_18889_ _11311_ _11312_ VGND VGND VPWR VPWR _11313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_241_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20920_ _02465_ _02688_ _02689_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__and3_1
XFILLER_0_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer13 net194 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
Xrebuffer24 _07059_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__buf_4
Xrebuffer35 net216 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_1
Xrebuffer46 _02827_ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_1
Xrebuffer57 _11691_ VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__buf_6
XFILLER_0_117_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20851_ _02517_ _02616_ _02623_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__a21o_1
Xrebuffer68 _01501_ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer79 _01416_ VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__clkbuf_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23570_ clknet_leaf_104_clk net738 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20782_ _02556_ _02557_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22521_ _04200_ _04201_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22452_ _03713_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21403_ top_inst.grid_inst.data_path_wires\[17\]\[3\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22383_ top_inst.grid_inst.data_path_wires\[18\]\[5\] _03713_ VGND VGND VPWR VPWR
+ _04068_ sky130_fd_sc_hd__and2b_1
XFILLER_0_33_959 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24122_ clknet_leaf_12_clk _00655_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_21334_ _03024_ _03063_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__nor2_1
XFILLER_0_206_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_1182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24053_ clknet_leaf_34_clk _00586_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold540 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[31\] VGND
+ VGND VPWR VPWR net722 sky130_fd_sc_hd__dlygate4sd3_1
X_21265_ _03002_ _03003_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold551 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[15\] VGND
+ VGND VPWR VPWR net733 sky130_fd_sc_hd__dlygate4sd3_1
X_23004_ top_inst.skew_buff_inst.row\[0\].output_reg\[3\] _04583_ VGND VGND VPWR VPWR
+ _04594_ sky130_fd_sc_hd__or2_1
Xhold562 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[1\] VGND
+ VGND VPWR VPWR net744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 top_inst.axis_out_inst.out_buff_data\[7\] VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__dlygate4sd3_1
X_20216_ _02013_ _11689_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__or2_1
XFILLER_0_229_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold584 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[2\] VGND VGND
+ VPWR VPWR net766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 top_inst.deskew_buff_inst.col_input\[121\] VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__dlygate4sd3_1
X_21196_ _02923_ _02917_ _02935_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_15__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_4_15__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_229_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20147_ _01956_ _01957_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__xor2_1
XFILLER_0_141_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20078_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[27\] _01764_ VGND
+ VGND VPWR VPWR _01892_ sky130_fd_sc_hd__xnor2_1
XTAP_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23906_ clknet_leaf_37_clk _00439_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ _04876_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__buf_2
XTAP_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _04876_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__clkbuf_2
XTAP_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23837_ clknet_leaf_92_clk _00370_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14570_ _07258_ _07259_ _07260_ VGND VGND VPWR VPWR _07262_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23768_ clknet_leaf_66_clk _00301_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11782_ top_inst.axis_out_inst.out_buff_data\[70\] _04890_ VGND VGND VPWR VPWR _04891_
+ sky130_fd_sc_hd__or2_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13521_ _06190_ _06188_ _06202_ _06200_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__and4_1
X_22719_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[24\] _04215_ _04216_
+ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23699_ clknet_leaf_124_clk _00232_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16240_ _08791_ _08822_ _08823_ VGND VGND VPWR VPWR _08824_ sky130_fd_sc_hd__and3_1
X_13452_ _06210_ _05773_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__or2_1
XFILLER_0_193_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12403_ net319 _05243_ _05244_ _05234_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16171_ _08756_ _08725_ _08734_ _08733_ _08732_ VGND VGND VPWR VPWR _08757_ sky130_fd_sc_hd__o32ai_4
X_13383_ _06146_ _06155_ VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15122_ _07769_ _07770_ _07741_ _07742_ VGND VGND VPWR VPWR _07772_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12334_ net863 _05204_ _05205_ _05195_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19930_ _01673_ _01694_ _01750_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__and3_1
X_15053_ _07703_ _07704_ VGND VGND VPWR VPWR _07705_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12265_ net650 _05156_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__or2_1
XFILLER_0_181_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14004_ _06714_ _06721_ VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19861_ _01527_ _01683_ _01684_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__nand3b_1
X_12196_ top_inst.axis_out_inst.out_buff_data\[25\] _05115_ VGND VGND VPWR VPWR _05126_
+ sky130_fd_sc_hd__or2_1
Xoutput60 net60 VGND VGND VPWR VPWR output_tdata[11] sky130_fd_sc_hd__clkbuf_4
Xoutput71 net71 VGND VGND VPWR VPWR output_tdata[14] sky130_fd_sc_hd__clkbuf_4
Xoutput82 net82 VGND VGND VPWR VPWR output_tdata[24] sky130_fd_sc_hd__clkbuf_4
X_18812_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[4\] _11210_ _11211_
+ VGND VGND VPWR VPWR _11238_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_128_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput93 net93 VGND VGND VPWR VPWR output_tdata[34] sky130_fd_sc_hd__clkbuf_4
X_19792_ _01617_ _01618_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__and2_1
XTAP_6061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18743_ _11170_ _11171_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[1\]
+ VGND VGND VPWR VPWR _11173_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15955_ _08484_ _08564_ VGND VGND VPWR VPWR _08565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_223_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14906_ _07579_ _07588_ VGND VGND VPWR VPWR _07589_ sky130_fd_sc_hd__xnor2_1
XTAP_5393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18674_ net948 _11116_ net167 VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__o21a_1
XTAP_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15886_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[10\] _08452_ _08373_
+ VGND VGND VPWR VPWR _08498_ sky130_fd_sc_hd__a21o_1
XTAP_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17625_ top_inst.grid_inst.data_path_wires\[11\]\[5\] top_inst.grid_inst.data_path_wires\[11\]\[4\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _10137_ sky130_fd_sc_hd__nand4_1
X_14837_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[14\] _07364_ VGND
+ VGND VPWR VPWR _07522_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_203_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17556_ _05732_ VGND VGND VPWR VPWR _10071_ sky130_fd_sc_hd__buf_4
X_14768_ _07449_ _07454_ VGND VGND VPWR VPWR _07455_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16507_ _09082_ _09083_ VGND VGND VPWR VPWR _09084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13719_ _06462_ _06449_ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__and2b_1
XFILLER_0_184_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17487_ _10014_ _10019_ _10020_ VGND VGND VPWR VPWR _10021_ sky130_fd_sc_hd__a21o_1
X_14699_ _07372_ _07373_ _07386_ VGND VGND VPWR VPWR _07388_ sky130_fd_sc_hd__nand3_1
XFILLER_0_73_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19226_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[15\] _10616_ _11640_
+ _11641_ VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16438_ _09015_ _09016_ VGND VGND VPWR VPWR _09017_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19157_ _11572_ _11574_ VGND VGND VPWR VPWR _11575_ sky130_fd_sc_hd__xor2_1
X_16369_ _08905_ _08907_ VGND VGND VPWR VPWR _08950_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18108_ _10591_ VGND VGND VPWR VPWR _10592_ sky130_fd_sc_hd__clkbuf_4
X_19088_ _11494_ _11468_ VGND VGND VPWR VPWR _11507_ sky130_fd_sc_hd__or2b_1
XFILLER_0_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18039_ _05309_ VGND VGND VPWR VPWR _10541_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21050_ _02643_ _02792_ _02503_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_61_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20001_ net1094 _01202_ _01817_ _01818_ _11228_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__o221a_1
XFILLER_0_226_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21952_ _03597_ _03616_ _03453_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_1103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20903_ _02004_ _02018_ _02438_ _02227_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__a31oi_4
X_21883_ _03574_ _03578_ _03600_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__nand3_1
XFILLER_0_94_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23622_ clknet_leaf_102_clk net263 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20834_ _02583_ _02584_ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23553_ clknet_leaf_105_clk _00086_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20765_ _02535_ _02541_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22504_ _04153_ _04184_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23484_ clknet_leaf_137_clk _00017_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[74\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20696_ _02472_ _02474_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22435_ _04115_ _04117_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22366_ _03926_ _03972_ _04050_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__and3_1
XFILLER_0_241_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24105_ clknet_leaf_15_clk _00638_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21317_ _03009_ _03054_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22297_ top_inst.grid_inst.data_path_wires\[18\]\[6\] top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[18\]\[7\]
+ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__a22o_1
X_24036_ clknet_leaf_41_clk _00569_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_12050_ net274 _05036_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold370 _00099_ VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__dlygate4sd3_1
X_21248_ _02963_ _02987_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__nand2_1
XFILLER_0_241_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold381 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[11\] VGND
+ VGND VPWR VPWR net563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold392 _00151_ VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__dlygate4sd3_1
X_21179_ _01819_ _02920_ _02921_ _02909_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15740_ _08352_ _08354_ VGND VGND VPWR VPWR _08355_ sky130_fd_sc_hd__nor2_2
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _05748_ _05735_ _05749_ _05743_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__o211a_1
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11903_ net430 _04951_ _04959_ _04955_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _08285_ _08286_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[6\]
+ VGND VGND VPWR VPWR _08288_ sky130_fd_sc_hd__a21oi_1
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _05687_ _05688_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__nor2_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17410_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[26\] _09496_ _09932_
+ _09948_ VGND VGND VPWR VPWR _09949_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14622_ _05632_ _07312_ VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _10606_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[5\] VGND
+ VGND VPWR VPWR _10855_ sky130_fd_sc_hd__nand2_1
X_11834_ net944 _04912_ _04920_ _04916_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__o211a_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17341_ _09867_ _09882_ VGND VGND VPWR VPWR _09883_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14553_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[5\] _07069_ _07243_
+ _07244_ VGND VGND VPWR VPWR _07245_ sky130_fd_sc_hd__nand4_1
X_11765_ top_inst.axis_out_inst.out_buff_data\[127\] _04877_ VGND VGND VPWR VPWR _04881_
+ sky130_fd_sc_hd__or2_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _06251_ _06254_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17272_ _09816_ _09809_ VGND VGND VPWR VPWR _09817_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14484_ _07169_ _07170_ _07177_ VGND VGND VPWR VPWR _07178_ sky130_fd_sc_hd__and3_1
X_19011_ _11147_ _11154_ _11396_ _11397_ VGND VGND VPWR VPWR _11432_ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16223_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[5\] _08773_ _08774_
+ VGND VGND VPWR VPWR _08807_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13435_ _06198_ _05262_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer4 _05265_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_181_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13366_ _05311_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__clkbuf_16
X_16154_ _05887_ _08738_ _08739_ _08740_ VGND VGND VPWR VPWR _08741_ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_942 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15105_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[5\] _07722_ _07723_
+ VGND VGND VPWR VPWR _07755_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_140_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12317_ _05142_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_239_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13297_ _06025_ _06072_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__xnor2_1
X_16085_ _08682_ VGND VGND VPWR VPWR _08683_ sky130_fd_sc_hd__buf_2
XFILLER_0_107_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15036_ _07688_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__clkbuf_1
X_12248_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[14\] _05156_
+ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__or2_1
X_19913_ net907 _10616_ _01734_ _11714_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19844_ _01656_ _01668_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__xor2_1
XFILLER_0_43_1084 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12179_ net485 _05115_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__or2_1
XFILLER_0_208_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19775_ _01528_ _01601_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__xor2_1
X_16987_ _09503_ _09502_ VGND VGND VPWR VPWR _09541_ sky130_fd_sc_hd__and2b_1
XFILLER_0_208_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18726_ _11140_ _10607_ _11159_ _11160_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15938_ _08509_ _08548_ VGND VGND VPWR VPWR _08549_ sky130_fd_sc_hd__xor2_2
XFILLER_0_223_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18657_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[16\] _10639_ VGND
+ VGND VPWR VPWR _11115_ sky130_fd_sc_hd__or2_1
X_15869_ _08443_ _08447_ VGND VGND VPWR VPWR _08481_ sky130_fd_sc_hd__nand2_1
XFILLER_0_203_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17608_ _10118_ _10120_ VGND VGND VPWR VPWR _10121_ sky130_fd_sc_hd__xor2_2
XFILLER_0_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18588_ _10969_ _11047_ VGND VGND VPWR VPWR _11048_ sky130_fd_sc_hd__xor2_1
XFILLER_0_175_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17539_ _10056_ _10057_ VGND VGND VPWR VPWR _10058_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20550_ _02330_ _02332_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_184_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19209_ _11514_ _11623_ VGND VGND VPWR VPWR _11625_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20481_ _02264_ _02265_ _05732_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22220_ _03709_ _03684_ _03869_ _03908_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22151_ _03840_ _03841_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21102_ _02862_ _11133_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__or2_1
XFILLER_0_199_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1054 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22082_ _03773_ _03774_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__nor2_1
XFILLER_0_199_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21033_ _02771_ _02772_ _02769_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__o21a_1
XFILLER_0_196_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_242_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22984_ net969 _04575_ _04582_ _04577_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21935_ _03618_ _03617_ _03633_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21866_ _03534_ _03582_ _03585_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23605_ clknet_leaf_104_clk _00138_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_20817_ _02590_ _02591_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24585_ clknet_leaf_20_clk _01118_ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dfxtp_4
X_21797_ _03499_ _03518_ _03512_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__nand3_1
XFILLER_0_194_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23536_ clknet_leaf_139_clk _00069_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_20748_ _02496_ _02524_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23467_ clknet_leaf_31_clk net778 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[121\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20679_ _02429_ _02434_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13220_ _05995_ _05997_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__xnor2_1
X_22418_ _04100_ _04101_ VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_190_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23398_ net842 _04655_ _04818_ _04819_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__o211a_1
X_13151_ _05744_ _05768_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22349_ _03991_ _03993_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12102_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[16\] _05063_
+ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__or2_1
XFILLER_0_221_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13082_ _05853_ _05862_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_237_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24019_ clknet_leaf_54_clk _00552_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_16910_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[3\]
+ _09210_ VGND VGND VPWR VPWR _09466_ sky130_fd_sc_hd__and3_1
X_12033_ net268 _05031_ _05033_ _05022_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17890_ _10350_ _10351_ _10395_ VGND VGND VPWR VPWR _10396_ sky130_fd_sc_hd__o21a_1
XFILLER_0_218_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16841_ _09393_ _09394_ _09395_ VGND VGND VPWR VPWR _09399_ sky130_fd_sc_hd__or3_1
XFILLER_0_232_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19560_ _01350_ _01356_ _01391_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16772_ _09324_ _09329_ _09330_ VGND VGND VPWR VPWR _09331_ sky130_fd_sc_hd__nand3_2
X_13984_ _06364_ _06702_ VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__and2_1
XFILLER_0_232_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18511_ _10971_ _10972_ VGND VGND VPWR VPWR _10973_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15723_ _08297_ _08298_ VGND VGND VPWR VPWR _08339_ sky130_fd_sc_hd__nor2_1
X_12935_ _05734_ _05735_ _05737_ _05308_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__o211a_1
X_19491_ _01306_ _01323_ _01324_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__nand3_1
XFILLER_0_125_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18442_ _10904_ _10905_ VGND VGND VPWR VPWR _10906_ sky130_fd_sc_hd__or2_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _08257_ _08259_ VGND VGND VPWR VPWR _08271_ sky130_fd_sc_hd__nand2_1
X_12866_ _05302_ _05305_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _07294_ _07295_ VGND VGND VPWR VPWR _07296_ sky130_fd_sc_hd__nand2_2
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11817_ top_inst.axis_out_inst.out_buff_data\[86\] _04903_ VGND VGND VPWR VPWR _04910_
+ sky130_fd_sc_hd__or2_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18373_ _10789_ _10795_ VGND VGND VPWR VPWR _10838_ sky130_fd_sc_hd__or2b_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15585_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[3\] _08203_ _08204_
+ VGND VGND VPWR VPWR _08205_ sky130_fd_sc_hd__and3_1
XFILLER_0_205_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12797_ _05293_ _05288_ _05305_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__and3_1
XFILLER_0_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _09866_ VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__clkbuf_1
X_14536_ _07200_ _07202_ VGND VGND VPWR VPWR _07228_ sky130_fd_sc_hd__nand2_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11748_ _04869_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__buf_8
XFILLER_0_83_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17255_ _09789_ _09800_ VGND VGND VPWR VPWR _09801_ sky130_fd_sc_hd__xnor2_1
X_14467_ _07113_ _07132_ _07154_ _07155_ VGND VGND VPWR VPWR _07161_ sky130_fd_sc_hd__and4b_1
XFILLER_0_183_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16206_ _08790_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13418_ _06186_ _05262_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__or2_1
X_17186_ _09733_ _09734_ _09726_ VGND VGND VPWR VPWR _09735_ sky130_fd_sc_hd__a21oi_1
X_14398_ _07066_ _07061_ _07065_ _07062_ VGND VGND VPWR VPWR _07096_ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16137_ _08688_ _08664_ _08661_ _08690_ VGND VGND VPWR VPWR _08724_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13349_ _06054_ _06122_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16068_ _08143_ _08663_ _08670_ _08666_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15019_ _07669_ _07671_ VGND VGND VPWR VPWR _07672_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_242_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19827_ _01518_ _01649_ _01651_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_235_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19758_ _01582_ _01583_ _01584_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_189_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18709_ _10595_ _11142_ _11148_ _11137_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__o211a_1
X_19689_ _01345_ _01514_ _01515_ _01517_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__o211a_4
XFILLER_0_211_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21720_ _03423_ _03426_ _03425_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_177_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21651_ _03246_ _03378_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__and2_1
XFILLER_0_231_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20602_ net795 _01735_ _02383_ _02035_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__o211a_1
X_24370_ clknet_leaf_40_clk net579 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[3\].output_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21582_ _03301_ _03280_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__or2b_1
XFILLER_0_117_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23321_ net152 _04766_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20533_ _01995_ _02227_ _02284_ _02285_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_172_661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23252_ net119 _04727_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20464_ _02246_ _02247_ _02240_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__a21o_1
XFILLER_0_171_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22203_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[1\] _03697_ top_inst.grid_inst.data_path_wires\[18\]\[7\]
+ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_30_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23183_ net86 _04687_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20395_ _01986_ _02178_ _02179_ _02180_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22134_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[18\]\[3\]
+ top_inst.grid_inst.data_path_wires\[18\]\[2\] _03707_ VGND VGND VPWR VPWR _03825_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_242_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22065_ top_inst.grid_inst.data_path_wires\[18\]\[3\] top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[1\]
+ _03697_ top_inst.grid_inst.data_path_wires\[18\]\[4\] VGND VGND VPWR VPWR _03758_
+ sky130_fd_sc_hd__a22o_1
XTAP_6649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21016_ _02782_ VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__clkbuf_1
XTAP_5937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_214_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22967_ top_inst.skew_buff_inst.row\[1\].output_reg\[3\] _04570_ VGND VGND VPWR VPWR
+ _04573_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12720_ _05527_ _05529_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21918_ _03628_ _03634_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__or2b_1
XFILLER_0_70_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22898_ net746 _04522_ _04533_ _04524_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12651_ _05280_ _05301_ _05305_ _05273_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24637_ clknet_leaf_26_clk _01170_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[113\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21849_ net524 _02638_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12582_ _05342_ _05355_ _05370_ _05395_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__o31a_1
X_15370_ _07973_ _07972_ VGND VGND VPWR VPWR _08014_ sky130_fd_sc_hd__or2b_1
XFILLER_0_108_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24568_ clknet_leaf_134_clk _01101_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14321_ _07027_ _07028_ _07029_ VGND VGND VPWR VPWR _07030_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_147_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23519_ clknet_leaf_138_clk net819 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1002 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24499_ clknet_leaf_128_clk _01032_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_184_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17040_ _09591_ _09592_ VGND VGND VPWR VPWR _09593_ sky130_fd_sc_hd__xor2_1
XFILLER_0_191_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14252_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[7\] VGND VGND
+ VPWR VPWR _06963_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13203_ _05979_ _05980_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__xor2_1
XFILLER_0_81_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1068 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14183_ _06850_ _06853_ _06851_ VGND VGND VPWR VPWR _06896_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_0_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13134_ _05911_ _05913_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18991_ _11393_ _11412_ VGND VGND VPWR VPWR _11413_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_238_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _05352_ _05846_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__and2_1
X_17942_ _04868_ VGND VGND VPWR VPWR _10447_ sky130_fd_sc_hd__buf_4
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12016_ net631 _05018_ _05024_ _05022_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17873_ _10035_ _10378_ _10059_ _10056_ VGND VGND VPWR VPWR _10379_ sky130_fd_sc_hd__and4_1
XFILLER_0_217_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16824_ _09338_ _09380_ _09381_ VGND VGND VPWR VPWR _09382_ sky130_fd_sc_hd__nand3_1
XFILLER_0_178_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19612_ _11697_ _01441_ _01442_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_233_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19543_ _01357_ _01374_ _01375_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16755_ _09278_ _09280_ VGND VGND VPWR VPWR _09315_ sky130_fd_sc_hd__nand2_1
X_13967_ top_inst.grid_inst.data_path_wires\[3\]\[4\] top_inst.grid_inst.data_path_wires\[3\]\[3\]
+ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[1\] top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__nand4_1
XFILLER_0_159_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15706_ _08316_ _08321_ VGND VGND VPWR VPWR _08322_ sky130_fd_sc_hd__xnor2_1
X_12918_ _05655_ _05712_ _05721_ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__a21o_1
X_19474_ _11688_ _11700_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16686_ _09194_ _09197_ _09202_ _09188_ VGND VGND VPWR VPWR _09248_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_232_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13898_ _06193_ _06192_ _06631_ _06446_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18425_ _10885_ _10888_ VGND VGND VPWR VPWR _10889_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15637_ _08248_ _08254_ VGND VGND VPWR VPWR _08255_ sky130_fd_sc_hd__xnor2_2
X_12849_ _05654_ _05605_ _05606_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__or3_1
XFILLER_0_115_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_232_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18356_ _10818_ _10821_ VGND VGND VPWR VPWR _10822_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_174_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15568_ _08187_ _08188_ VGND VGND VPWR VPWR _08189_ sky130_fd_sc_hd__xnor2_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17307_ _09822_ _09847_ VGND VGND VPWR VPWR _09850_ sky130_fd_sc_hd__and2b_1
XFILLER_0_127_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14519_ _07198_ _07199_ _07209_ _07210_ VGND VGND VPWR VPWR _07212_ sky130_fd_sc_hd__a22o_1
XFILLER_0_173_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18287_ _10729_ _10730_ VGND VGND VPWR VPWR _10754_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15499_ top_inst.grid_inst.data_path_wires\[7\]\[1\] VGND VGND VPWR VPWR _08137_
+ sky130_fd_sc_hd__buf_4
XFILLER_0_182_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17238_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[18\] _09496_ _09783_
+ _09784_ VGND VGND VPWR VPWR _09785_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_834 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold903 top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[13\] VGND VGND
+ VPWR VPWR net1085 sky130_fd_sc_hd__dlygate4sd3_1
X_17169_ _09690_ _09715_ VGND VGND VPWR VPWR _09718_ sky130_fd_sc_hd__nand2_1
Xhold914 top_inst.deskew_buff_inst.col_input\[17\] VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold925 top_inst.axis_out_inst.out_buff_data\[99\] VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20180_ _01987_ _10033_ _01988_ _01840_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23870_ clknet_leaf_78_clk _00403_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22821_ _04364_ _04459_ _04461_ _04486_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__a211o_1
XFILLER_0_212_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22752_ _05312_ _04409_ _04420_ _04421_ _04422_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__a41o_1
XFILLER_0_17_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21703_ _03428_ _03429_ VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__xnor2_2
X_22683_ _04334_ _04356_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_133_1262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24422_ clknet_leaf_56_clk _00955_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21634_ _03314_ _03334_ _03363_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_136_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24353_ clknet_leaf_26_clk _00886_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[112\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21565_ _03210_ _03260_ _03296_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23304_ net144 _04766_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__or2_1
X_20516_ _02297_ _02298_ _02282_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__a21o_1
X_24284_ clknet_leaf_10_clk _00817_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21496_ _03227_ _03229_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__xor2_2
XFILLER_0_144_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23235_ net111 _04727_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__or2_1
X_20447_ _01990_ _02229_ _02230_ _02231_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__o22a_1
XFILLER_0_209_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23166_ net382 _04685_ _04688_ _04675_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20378_ _02162_ _02163_ _02120_ _02122_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__o211a_1
XTAP_6402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22117_ _03795_ _03797_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23097_ net605 _05323_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_237_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22048_ _03739_ _03741_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__nand2_1
XFILLER_0_238_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14870_ _07553_ _07554_ _06682_ VGND VGND VPWR VPWR _07555_ sky130_fd_sc_hd__a21o_1
XTAP_5789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13821_ _06526_ _06530_ _06561_ VGND VGND VPWR VPWR _06563_ sky130_fd_sc_hd__or3_1
XFILLER_0_230_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23999_ clknet_leaf_81_clk net1069 VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_106_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_214_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16540_ _09080_ _09048_ _09090_ VGND VGND VPWR VPWR _09116_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13752_ _06494_ _06495_ VGND VGND VPWR VPWR _06496_ sky130_fd_sc_hd__nor2_2
XFILLER_0_98_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12703_ _05512_ _05513_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__and2_1
XFILLER_0_168_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16471_ _09007_ _09047_ VGND VGND VPWR VPWR _09049_ sky130_fd_sc_hd__or2_1
X_13683_ _06428_ _06378_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1069 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18210_ _10678_ _10679_ VGND VGND VPWR VPWR _10680_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15422_ _08061_ _08063_ _08064_ VGND VGND VPWR VPWR _08065_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12634_ _05413_ _05414_ _05420_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__and3_1
X_19190_ _11588_ _11606_ VGND VGND VPWR VPWR _11607_ sky130_fd_sc_hd__or2b_1
XFILLER_0_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18141_ _10595_ _10607_ _10615_ _10594_ VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15353_ _07995_ _07996_ VGND VGND VPWR VPWR _07997_ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12565_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[3\]
+ _05279_ _05282_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__nand4_1
XFILLER_0_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14304_ _07012_ _07013_ VGND VGND VPWR VPWR _07014_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18072_ _10565_ _10571_ VGND VGND VPWR VPWR _10572_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15284_ _07923_ _07929_ VGND VGND VPWR VPWR _07930_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12496_ _05310_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__buf_6
XFILLER_0_41_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17023_ _09540_ _09535_ _09576_ VGND VGND VPWR VPWR _09577_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14235_ _06945_ _06946_ VGND VGND VPWR VPWR _06947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14166_ _06836_ _06838_ _06879_ VGND VGND VPWR VPWR _06880_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1032 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13117_ top_inst.grid_inst.data_path_wires\[1\]\[5\] _05761_ _05895_ _05896_ VGND
+ VGND VPWR VPWR _05897_ sky130_fd_sc_hd__a22o_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14097_ _06772_ _06773_ VGND VGND VPWR VPWR _06812_ sky130_fd_sc_hd__nor2_1
X_18974_ top_inst.grid_inst.data_path_wires\[13\]\[5\] _11158_ _11156_ top_inst.grid_inst.data_path_wires\[13\]\[6\]
+ VGND VGND VPWR VPWR _11396_ sky130_fd_sc_hd__a22o_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _05746_ _05744_ _05759_ _05757_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__and4_1
X_17925_ _10428_ _10429_ VGND VGND VPWR VPWR _10430_ sky130_fd_sc_hd__nand2_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17856_ net1083 _09494_ VGND VGND VPWR VPWR _10363_ sky130_fd_sc_hd__or2_1
XFILLER_0_179_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16807_ _09193_ _09188_ _09215_ net219 VGND VGND VPWR VPWR _09365_ sky130_fd_sc_hd__nand4_1
XFILLER_0_89_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17787_ _10292_ _10294_ VGND VGND VPWR VPWR _10295_ sky130_fd_sc_hd__and2_1
X_14999_ _07652_ _07653_ _06682_ VGND VGND VPWR VPWR _07654_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16738_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[5\] _09296_ _09297_
+ VGND VGND VPWR VPWR _09298_ sky130_fd_sc_hd__and3_1
XFILLER_0_163_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19526_ _11697_ _11696_ _11700_ _11693_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_92_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19457_ _01195_ _01221_ _01222_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__and3_1
X_16669_ _09198_ _09187_ VGND VGND VPWR VPWR _09232_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18408_ _10788_ _10817_ _10872_ VGND VGND VPWR VPWR _10873_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19388_ _01223_ _01224_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18339_ _10803_ _10804_ VGND VGND VPWR VPWR _10805_ sky130_fd_sc_hd__and2b_1
XFILLER_0_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21350_ _02875_ _02887_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20301_ _01987_ _02016_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[4\]
+ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_163_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold700 _00963_ VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__dlygate4sd3_1
X_21281_ _02997_ _03018_ _03019_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__and3_1
Xhold711 top_inst.deskew_buff_inst.col_input\[106\] VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold722 _00974_ VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__dlygate4sd3_1
X_23020_ net1 _04601_ _04604_ _04590_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold733 _00091_ VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__dlygate4sd3_1
X_20232_ _01987_ _02007_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__a21oi_1
Xhold744 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[14\] VGND
+ VGND VPWR VPWR net926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 _00902_ VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold766 top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[18\] VGND VGND
+ VPWR VPWR net948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[19\] VGND VGND
+ VPWR VPWR net959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20163_ _01951_ _01955_ _01953_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__a21oi_1
Xhold788 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[6\] VGND
+ VGND VPWR VPWR net970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold799 top_inst.deskew_buff_inst.col_input\[27\] VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__buf_1
XFILLER_0_25_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20094_ _01882_ _01885_ _01906_ _10957_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__a31o_1
XFILLER_0_239_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23922_ clknet_leaf_77_clk _00455_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23853_ clknet_leaf_68_clk _00386_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22804_ _04467_ _04471_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23784_ clknet_leaf_65_clk _00317_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_20996_ _02715_ _02760_ _02762_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__o21a_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22735_ net777 _05317_ _04405_ _04406_ _09806_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__o221a_1
XFILLER_0_32_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22666_ top_inst.deskew_buff_inst.col_input\[118\] _05731_ _04326_ _04340_ VGND VGND
+ VPWR VPWR _04341_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24405_ clknet_leaf_39_clk net417 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].output_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21617_ _03305_ _03338_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22597_ _04273_ _04274_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12350_ net747 _05204_ _05214_ _05208_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__o211a_1
X_24336_ clknet_leaf_5_clk _00869_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_21548_ _03279_ _03247_ _03249_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_244_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_244_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12281_ net695 _05169_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24267_ clknet_leaf_101_clk _00800_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_21479_ top_inst.grid_inst.data_path_wires\[17\]\[5\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14020_ _06714_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__inv_2
X_23218_ net613 _04713_ _04718_ _04717_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24198_ clknet_leaf_116_clk _00731_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23149_ net71 _04672_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15971_ _08531_ _08536_ _08534_ VGND VGND VPWR VPWR _08581_ sky130_fd_sc_hd__a21o_1
XTAP_6265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17710_ _10194_ _10219_ VGND VGND VPWR VPWR _10220_ sky130_fd_sc_hd__xnor2_1
XTAP_6298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14922_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[21\] _07595_ VGND
+ VGND VPWR VPWR _07600_ sky130_fd_sc_hd__and2_1
XTAP_5553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18690_ top_inst.grid_inst.data_path_wires\[13\]\[2\] VGND VGND VPWR VPWR _11135_
+ sky130_fd_sc_hd__clkbuf_4
XTAP_5575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold82 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[23\] VGND
+ VGND VPWR VPWR net264 sky130_fd_sc_hd__dlygate4sd3_1
X_17641_ _09661_ _10152_ VGND VGND VPWR VPWR _10153_ sky130_fd_sc_hd__and2_1
X_14853_ _07526_ _07537_ VGND VGND VPWR VPWR _07538_ sky130_fd_sc_hd__xor2_1
XFILLER_0_216_1112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold93 _00161_ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _06467_ _06514_ _06512_ VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__a21oi_1
X_17572_ _10076_ _10077_ VGND VGND VPWR VPWR _10086_ sky130_fd_sc_hd__or2b_1
XFILLER_0_231_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14784_ _07470_ VGND VGND VPWR VPWR _07471_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11996_ net556 _05010_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__or2_1
X_19311_ _11707_ VGND VGND VPWR VPWR _11708_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16523_ _09091_ _09092_ _09098_ VGND VGND VPWR VPWR _09100_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13735_ _06447_ _06443_ _06479_ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__a21o_1
XFILLER_0_202_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19242_ _11630_ _11631_ _11656_ VGND VGND VPWR VPWR _11657_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16454_ _09001_ _09002_ _09031_ VGND VGND VPWR VPWR _09033_ sky130_fd_sc_hd__or3_1
XFILLER_0_112_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13666_ _06188_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[6\] _06410_
+ VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15405_ _08043_ _08047_ VGND VGND VPWR VPWR _08048_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12617_ _05428_ _05429_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__or2_1
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19173_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[14\] _11469_ VGND
+ VGND VPWR VPWR _11590_ sky130_fd_sc_hd__and2_1
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16385_ _08922_ _08924_ _08921_ VGND VGND VPWR VPWR _08965_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_213_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13597_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[7\] _06342_ _06344_
+ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18124_ _10581_ _10046_ _10603_ _10594_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15336_ _07978_ _07980_ VGND VGND VPWR VPWR _07981_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12548_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[3\]
+ _05271_ _05278_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18055_ _10554_ _10555_ VGND VGND VPWR VPWR _10556_ sky130_fd_sc_hd__nand2_1
X_15267_ _07911_ _07912_ VGND VGND VPWR VPWR _07913_ sky130_fd_sc_hd__xnor2_1
X_12479_ top_inst.skew_buff_inst.row\[0\].output_reg\[6\] top_inst.axis_in_inst.inbuf_bus\[6\]
+ _05267_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__mux2_1
XANTENNA_2 _05044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17006_ _09557_ _09558_ _09559_ VGND VGND VPWR VPWR _09560_ sky130_fd_sc_hd__and3_1
X_14218_ _06928_ _06929_ VGND VGND VPWR VPWR _06930_ sky130_fd_sc_hd__xnor2_1
X_15198_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[8\] _07845_ VGND
+ VGND VPWR VPWR _07846_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14149_ _06813_ VGND VGND VPWR VPWR _06863_ sky130_fd_sc_hd__inv_2
XFILLER_0_201_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18957_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[8\] _09496_ _11378_
+ _11379_ VGND VGND VPWR VPWR _11380_ sky130_fd_sc_hd__a22o_1
XFILLER_0_226_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17908_ _10412_ VGND VGND VPWR VPWR _10413_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18888_ _11143_ _11154_ _11309_ _11310_ VGND VGND VPWR VPWR _11312_ sky130_fd_sc_hd__nand4_1
XFILLER_0_94_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer14 _01458_ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_1
X_17839_ _10338_ _10345_ VGND VGND VPWR VPWR _10346_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_234_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer25 net206 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__buf_1
XFILLER_0_89_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer36 _01234_ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__buf_1
XFILLER_0_117_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer47 _01464_ VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__buf_2
X_20850_ _02518_ _02622_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__xnor2_1
Xrebuffer58 net239 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer69 net250 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19509_ top_inst.deskew_buff_inst.col_input\[7\] _01342_ _08307_ VGND VGND VPWR VPWR
+ _01343_ sky130_fd_sc_hd__mux2_1
X_20781_ _02517_ _02548_ _02555_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__nand3_1
XFILLER_0_193_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22520_ _04137_ _04199_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22451_ _04025_ _04107_ _04133_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__a21o_1
XFILLER_0_228_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21402_ top_inst.grid_inst.data_path_wires\[17\]\[2\] _02897_ VGND VGND VPWR VPWR
+ _03138_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22382_ _03695_ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[5\] VGND
+ VGND VPWR VPWR _04067_ sky130_fd_sc_hd__and2_1
XFILLER_0_228_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24121_ clknet_leaf_13_clk _00654_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_21333_ _07057_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__buf_4
XFILLER_0_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold530 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[7\] VGND VGND
+ VPWR VPWR net712 sky130_fd_sc_hd__dlygate4sd3_1
X_24052_ clknet_leaf_34_clk _00585_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21264_ _03000_ _03001_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[6\]
+ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold541 top_inst.axis_out_inst.out_buff_data\[26\] VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[0\] VGND VGND
+ VPWR VPWR net734 sky130_fd_sc_hd__dlygate4sd3_1
X_23003_ net951 _04588_ _04593_ _04590_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold563 top_inst.deskew_buff_inst.col_input\[39\] VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__dlygate4sd3_1
X_20215_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[3\] VGND VGND
+ VPWR VPWR _02013_ sky130_fd_sc_hd__buf_4
Xhold574 top_inst.deskew_buff_inst.col_input\[28\] VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__dlygate4sd3_1
X_21195_ _02936_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold585 _00936_ VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 _00000_ VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1057 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_239_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20146_ _01783_ _01939_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_239_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20077_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[26\] _01761_ _01762_
+ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__a21o_2
XTAP_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23905_ clknet_leaf_54_clk _00438_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23836_ clknet_leaf_92_clk _00369_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11850_ net313 _04925_ _04928_ _04929_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23767_ clknet_leaf_66_clk _00300_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11781_ _04876_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__buf_2
XFILLER_0_67_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20979_ _02718_ _02746_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13520_ _06264_ _06269_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__xor2_2
X_22718_ _04388_ _04389_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__nand2_2
XFILLER_0_94_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23698_ clknet_leaf_124_clk _00231_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13451_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[4\] VGND VGND
+ VPWR VPWR _06210_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22649_ net260 _03528_ _04323_ _04324_ _09806_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__o221a_1
XFILLER_0_137_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12402_ top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[17\] _05235_
+ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16170_ _08724_ VGND VGND VPWR VPWR _08756_ sky130_fd_sc_hd__inv_2
X_13382_ _06099_ _06154_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15121_ _07741_ _07742_ _07769_ _07770_ VGND VGND VPWR VPWR _07771_ sky130_fd_sc_hd__a211o_1
XFILLER_0_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24319_ clknet_leaf_139_clk _00852_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[94\]
+ sky130_fd_sc_hd__dfxtp_1
X_12333_ net329 _05196_ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_1283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15052_ _07681_ _07684_ VGND VGND VPWR VPWR _07704_ sky130_fd_sc_hd__nand2_1
XFILLER_0_239_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12264_ net958 _05164_ _05165_ _05155_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14003_ _06715_ _06720_ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19860_ _01394_ _01524_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[17\]
+ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__a21o_1
X_12195_ net900 _05123_ _05125_ _05114_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput50 net50 VGND VGND VPWR VPWR output_tdata[110] sky130_fd_sc_hd__clkbuf_4
Xoutput61 net61 VGND VGND VPWR VPWR output_tdata[120] sky130_fd_sc_hd__clkbuf_4
X_18811_ _11231_ _11236_ VGND VGND VPWR VPWR _11237_ sky130_fd_sc_hd__xnor2_2
Xoutput72 net72 VGND VGND VPWR VPWR output_tdata[15] sky130_fd_sc_hd__clkbuf_4
XTAP_6040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput83 net83 VGND VGND VPWR VPWR output_tdata[25] sky130_fd_sc_hd__clkbuf_4
XTAP_6051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19791_ _01599_ _01616_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__or2_1
Xoutput94 net94 VGND VGND VPWR VPWR output_tdata[35] sky130_fd_sc_hd__clkbuf_4
XTAP_6062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18742_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[1\] _11170_ _11171_
+ VGND VGND VPWR VPWR _11172_ sky130_fd_sc_hd__nand3_1
X_15954_ _08562_ _08563_ VGND VGND VPWR VPWR _08564_ sky130_fd_sc_hd__xnor2_1
XTAP_6095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14905_ _07581_ _07587_ VGND VGND VPWR VPWR _07588_ sky130_fd_sc_hd__xnor2_1
XTAP_5383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18673_ net922 _11116_ net167 VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__o21a_1
XTAP_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15885_ _08495_ _08496_ VGND VGND VPWR VPWR _08497_ sky130_fd_sc_hd__or2b_1
XFILLER_0_215_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14836_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[13\] _07364_ _07280_
+ VGND VGND VPWR VPWR _07521_ sky130_fd_sc_hd__a21o_1
XFILLER_0_187_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17624_ top_inst.grid_inst.data_path_wires\[11\]\[4\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[0\] top_inst.grid_inst.data_path_wires\[11\]\[5\]
+ VGND VGND VPWR VPWR _10136_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_231_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ net867 _08183_ _10070_ _10049_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__o211a_1
X_14767_ _07452_ _07453_ VGND VGND VPWR VPWR _07454_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11979_ net720 _04990_ _05002_ _04995_ VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_1298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16506_ _08876_ _08677_ _09081_ VGND VGND VPWR VPWR _09083_ sky130_fd_sc_hd__nor3_1
X_13718_ _06449_ _06462_ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__and2b_1
X_17486_ _10014_ _10019_ _05316_ VGND VGND VPWR VPWR _10020_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14698_ _07372_ _07373_ _07386_ VGND VGND VPWR VPWR _07387_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16437_ _09007_ _09014_ VGND VGND VPWR VPWR _09016_ sky130_fd_sc_hd__or2_1
X_19225_ _10447_ VGND VGND VPWR VPWR _11641_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13649_ _06393_ _06395_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_229_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19156_ _11519_ _11534_ _11573_ VGND VGND VPWR VPWR _11574_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16368_ _08947_ _08948_ VGND VGND VPWR VPWR _08949_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18107_ top_inst.grid_inst.data_path_wires\[12\]\[6\] VGND VGND VPWR VPWR _10591_
+ sky130_fd_sc_hd__buf_2
X_15319_ _07962_ _07963_ VGND VGND VPWR VPWR _07964_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19087_ _11492_ _11493_ VGND VGND VPWR VPWR _11506_ sky130_fd_sc_hd__nand2_1
X_16299_ _08835_ _08836_ VGND VGND VPWR VPWR _08881_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_120_clk clknet_4_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18038_ _10520_ _10539_ VGND VGND VPWR VPWR _10540_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_998 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20000_ _01798_ _01816_ _09292_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_226_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19989_ _01783_ _01782_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_241_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21951_ _03629_ _03633_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__or2b_1
XFILLER_0_158_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20902_ _02671_ _02672_ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21882_ _03574_ _03578_ _03600_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23621_ clknet_leaf_102_clk net255 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_1327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20833_ _02605_ _02606_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23552_ clknet_leaf_129_clk _00085_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20764_ _02538_ _02539_ _02540_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__nor3_1
XFILLER_0_92_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22503_ _04152_ _04180_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23483_ clknet_leaf_134_clk net368 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[73\]
+ sky130_fd_sc_hd__dfxtp_1
X_20695_ _02469_ _02471_ _02473_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22434_ _04115_ _04117_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_208_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22365_ _04005_ _04046_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_111_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24104_ clknet_leaf_15_clk _00637_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_21316_ _03050_ _03053_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22296_ top_inst.grid_inst.data_path_wires\[18\]\[7\] top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _03983_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24035_ clknet_leaf_41_clk _00568_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21247_ _02984_ _02986_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__xor2_1
Xhold360 top_inst.deskew_buff_inst.col_input\[115\] VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 top_inst.axis_out_inst.out_buff_data\[48\] VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold382 top_inst.deskew_buff_inst.col_input\[124\] VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 top_inst.axis_out_inst.out_buff_data\[98\] VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21178_ net282 _02638_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_1131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20129_ _01939_ _01940_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_244_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_244_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_189_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _05739_ _05597_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__nand2_1
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11902_ top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[26\] _04956_
+ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__or2_1
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15670_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[6\] _08285_ _08286_
+ VGND VGND VPWR VPWR _08287_ sky130_fd_sc_hd__and3_1
X_12882_ _05685_ _05686_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[8\] _05634_ _07310_
+ _07311_ VGND VGND VPWR VPWR _07312_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_185_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23819_ clknet_leaf_93_clk _00352_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_11833_ net434 _04917_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__or2_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17340_ _09880_ _09881_ VGND VGND VPWR VPWR _09882_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14552_ _07241_ _07060_ _07064_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _07244_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_185_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ net471 _04860_ _04880_ _04875_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__o211a_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13503_ _06210_ _06252_ _06253_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__a21bo_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17271_ _09813_ _09815_ VGND VGND VPWR VPWR _09816_ sky130_fd_sc_hd__xor2_2
XFILLER_0_138_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14483_ _07175_ _07176_ VGND VGND VPWR VPWR _07177_ sky130_fd_sc_hd__nor2_1
XFILLER_0_193_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19010_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[9\] _11340_ _11387_
+ VGND VGND VPWR VPWR _11431_ sky130_fd_sc_hd__a21o_1
X_16222_ _08796_ _08805_ VGND VGND VPWR VPWR _08806_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13434_ top_inst.grid_inst.data_path_wires\[2\]\[7\] VGND VGND VPWR VPWR _06198_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer5 net186 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_1
X_16153_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[3\] _05730_ VGND
+ VGND VPWR VPWR _08740_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13365_ _06106_ _06109_ _06138_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_102_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_148_1389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15104_ _07717_ _07753_ VGND VGND VPWR VPWR _07754_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12316_ net875 _05191_ _05194_ _05195_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__o211a_1
X_16084_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[0\] VGND VGND
+ VPWR VPWR _08682_ sky130_fd_sc_hd__buf_2
XFILLER_0_122_954 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13296_ _06070_ _06071_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19912_ _01717_ _01732_ _01733_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__o21ai_2
X_15035_ _07117_ _07687_ VGND VGND VPWR VPWR _07688_ sky130_fd_sc_hd__and2_1
X_12247_ _05142_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_236_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19843_ _01657_ _01667_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__xnor2_1
X_12178_ net346 _05110_ _05116_ _05114_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_1096 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19774_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[14\] _01480_ VGND
+ VGND VPWR VPWR _01601_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16986_ _09497_ _09531_ VGND VGND VPWR VPWR _09540_ sky130_fd_sc_hd__or2_1
XFILLER_0_194_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18725_ _10447_ VGND VGND VPWR VPWR _11160_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_218_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15937_ _08546_ _08547_ VGND VGND VPWR VPWR _08548_ sky130_fd_sc_hd__nor2_1
XTAP_5191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15868_ _08442_ _08441_ VGND VGND VPWR VPWR _08480_ sky130_fd_sc_hd__or2b_1
X_18656_ _11097_ _11113_ VGND VGND VPWR VPWR _11114_ sky130_fd_sc_hd__xor2_1
XTAP_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_204_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14819_ _07493_ _07494_ _07504_ VGND VGND VPWR VPWR _07505_ sky130_fd_sc_hd__a21o_1
XFILLER_0_203_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17607_ _10095_ _10096_ _10119_ VGND VGND VPWR VPWR _10120_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_188_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15799_ _08360_ _08363_ _08364_ _08412_ _08357_ VGND VGND VPWR VPWR _08413_ sky130_fd_sc_hd__a32oi_4
X_18587_ _11045_ _11046_ VGND VGND VPWR VPWR _11047_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17538_ _05772_ VGND VGND VPWR VPWR _10057_ sky130_fd_sc_hd__buf_2
XFILLER_0_114_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17469_ _10001_ _09995_ _10004_ VGND VGND VPWR VPWR _10005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19208_ _11514_ _11623_ VGND VGND VPWR VPWR _11624_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_871 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20480_ _02221_ _02263_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19139_ _11524_ _11525_ _11527_ VGND VGND VPWR VPWR _11557_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22150_ _03838_ _03839_ _03806_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21101_ top_inst.grid_inst.data_path_wires\[17\]\[0\] VGND VGND VPWR VPWR _02862_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22081_ _03751_ _03753_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21032_ _02796_ _02797_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__and2_1
XFILLER_0_227_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_1030 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22983_ net772 _04570_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__or2_1
XFILLER_0_241_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21934_ _03637_ _03639_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__or2b_1
XFILLER_0_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21865_ _03561_ _03554_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__and2b_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23604_ clknet_leaf_104_clk _00137_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20816_ _02589_ _02569_ _02571_ _05406_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__a31o_1
X_24584_ clknet_leaf_141_clk _01117_ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dfxtp_1
X_21796_ _03499_ _03512_ _03518_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23535_ clknet_leaf_140_clk net562 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20747_ _02522_ _02523_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__nor2_1
XFILLER_0_231_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23466_ net441 _04859_ _04855_ _06180_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__o211a_1
X_20678_ _02449_ _02447_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__and2b_1
XFILLER_0_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22417_ top_inst.grid_inst.data_path_wires\[18\]\[6\] _03713_ VGND VGND VPWR VPWR
+ _04101_ sky130_fd_sc_hd__or2b_1
XFILLER_0_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_243_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23397_ _04869_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_162_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13150_ _05927_ _05928_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22348_ _04025_ _04033_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12101_ net587 _05071_ _05072_ _05062_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__o211a_1
X_13081_ _05856_ _05861_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22279_ _03964_ _03966_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24018_ clknet_leaf_54_clk _00551_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_12032_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[18\] _05023_
+ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__or2_1
Xhold190 _01157_ VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16840_ _09361_ _09396_ _09397_ VGND VGND VPWR VPWR _09398_ sky130_fd_sc_hd__or3b_1
XFILLER_0_219_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16771_ _09327_ _09328_ _09305_ _09306_ VGND VGND VPWR VPWR _09330_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_189_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13983_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[4\] _06700_ _06701_
+ VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_244_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15722_ _08335_ _08337_ VGND VGND VPWR VPWR _08338_ sky130_fd_sc_hd__xnor2_1
X_18510_ _10968_ _10970_ VGND VGND VPWR VPWR _10972_ sky130_fd_sc_hd__and2_1
X_12934_ _05736_ _05272_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__or2_1
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ _01321_ _01322_ _01307_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__a21o_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18441_ _10890_ _10891_ _10903_ VGND VGND VPWR VPWR _10905_ sky130_fd_sc_hd__and3_1
X_15653_ _08238_ _08256_ VGND VGND VPWR VPWR _08270_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12865_ _05643_ _05644_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.weight_reg\[5\] _07073_ _07291_
+ _07293_ VGND VGND VPWR VPWR _07295_ sky130_fd_sc_hd__a22o_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11816_ net908 _04898_ _04909_ _04902_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _10794_ _10790_ VGND VGND VPWR VPWR _10837_ sky130_fd_sc_hd__or2b_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _08143_ _08139_ _08157_ _08155_ VGND VGND VPWR VPWR _08204_ sky130_fd_sc_hd__nand4_1
X_12796_ _05293_ _05288_ _05306_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_200_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _09661_ _09865_ VGND VGND VPWR VPWR _09866_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14535_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[6\] _07192_ _07193_
+ VGND VGND VPWR VPWR _07227_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_141_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11747_ _04868_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__clkbuf_8
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17254_ _09798_ _09799_ VGND VGND VPWR VPWR _09800_ sky130_fd_sc_hd__xnor2_1
X_14466_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[5\] VGND VGND
+ VPWR VPWR _07160_ sky130_fd_sc_hd__inv_2
XFILLER_0_181_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16205_ _08197_ _08789_ VGND VGND VPWR VPWR _08790_ sky130_fd_sc_hd__and2_1
XFILLER_0_226_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13417_ top_inst.grid_inst.data_path_wires\[2\]\[2\] VGND VGND VPWR VPWR _06186_
+ sky130_fd_sc_hd__clkbuf_4
X_17185_ _09731_ _09732_ _09728_ VGND VGND VPWR VPWR _09734_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14397_ net1077 _06660_ _07095_ _07092_ VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16136_ _08714_ _08715_ VGND VGND VPWR VPWR _08723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13348_ _06120_ _06121_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16067_ _08669_ _08140_ VGND VGND VPWR VPWR _08670_ sky130_fd_sc_hd__or2_1
X_13279_ _06050_ _06054_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15018_ _07631_ _07670_ VGND VGND VPWR VPWR _07671_ sky130_fd_sc_hd__nand2_2
XFILLER_0_122_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_208_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19826_ _01594_ _01648_ _01650_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_208_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19757_ _01582_ _01583_ _01584_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__and3_1
XFILLER_0_159_1271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16969_ _09521_ _09522_ _09505_ VGND VGND VPWR VPWR _09524_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_224_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18708_ _11147_ _11133_ VGND VGND VPWR VPWR _11148_ sky130_fd_sc_hd__or2_1
X_19688_ _01516_ _01474_ _01510_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__a21o_1
XFILLER_0_231_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18639_ _11040_ _11070_ _11093_ _11096_ _11092_ VGND VGND VPWR VPWR _11097_ sky130_fd_sc_hd__a32o_1
XFILLER_0_231_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21650_ _03246_ _03378_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20601_ _02351_ _02381_ _02382_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21581_ _03300_ _03299_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__or2b_1
XFILLER_0_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23320_ net629 _04765_ _04775_ _04769_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__o211a_1
X_20532_ _02277_ _02279_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23251_ net821 _04726_ _04736_ _04730_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__o211a_1
X_20463_ _02240_ _02246_ _02247_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__nand3_1
XFILLER_0_162_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22202_ top_inst.grid_inst.data_path_wires\[18\]\[7\] top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _03891_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23182_ net768 _04685_ _04697_ _04691_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20394_ top_inst.grid_inst.data_path_wires\[16\]\[3\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[7\] VGND VGND VPWR VPWR
+ _02180_ sky130_fd_sc_hd__and3_1
XFILLER_0_242_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_203_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22133_ _03822_ _03823_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__nor2_1
XFILLER_0_203_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22064_ _03757_ VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21015_ _02135_ _02781_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22966_ net772 _04562_ _04572_ _04564_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21917_ _03629_ _03633_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22897_ net674 _04530_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_242_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12650_ _05284_ _05292_ _05418_ _05417_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__a31o_1
XFILLER_0_167_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24636_ clknet_leaf_25_clk net509 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[112\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21848_ _03549_ _03568_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__xor2_1
XFILLER_0_195_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12581_ _05345_ _05369_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__or2b_1
X_24567_ clknet_leaf_138_clk _01100_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_182_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21779_ _03501_ _03502_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14320_ _06963_ _06635_ _06966_ _06997_ VGND VGND VPWR VPWR _07029_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23518_ clknet_leaf_138_clk net840 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24498_ clknet_leaf_125_clk _01031_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_81_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1014 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14251_ _06932_ _06936_ VGND VGND VPWR VPWR _06962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23449_ top_inst.axis_out_inst.out_buff_data\[112\] _04835_ VGND VGND VPWR VPWR _04847_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_11_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13202_ _05753_ _05761_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__nand2_2
XFILLER_0_123_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14182_ _06893_ _06894_ VGND VGND VPWR VPWR _06895_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13133_ _05863_ _05871_ _05912_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18990_ _11410_ _11411_ VGND VGND VPWR VPWR _11412_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[5\] _05354_ _05844_
+ _05845_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__a22o_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ net1089 _09494_ VGND VGND VPWR VPWR _10446_ sky130_fd_sc_hd__or2_1
XFILLER_0_237_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12015_ net488 _05023_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__or2_1
X_17872_ top_inst.grid_inst.data_path_wires\[11\]\[4\] VGND VGND VPWR VPWR _10378_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_139_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19611_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[4\] _11704_ _11708_
+ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _01442_ sky130_fd_sc_hd__a22o_1
XFILLER_0_219_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16823_ _09378_ _09379_ _09376_ VGND VGND VPWR VPWR _09381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19542_ _01371_ _01372_ _01373_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__a21o_1
X_16754_ _09311_ _09312_ _09282_ VGND VGND VPWR VPWR _09314_ sky130_fd_sc_hd__o21a_1
X_13966_ _06672_ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__inv_2
XFILLER_0_232_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12917_ _05709_ _05711_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__and2b_1
X_15705_ _08319_ _08320_ VGND VGND VPWR VPWR _08321_ sky130_fd_sc_hd__nand2_1
X_16685_ _09237_ _09238_ VGND VGND VPWR VPWR _09247_ sky130_fd_sc_hd__nor2_1
X_19473_ _01272_ _01273_ _01276_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__and3_1
XFILLER_0_201_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13897_ _06630_ _06620_ VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18424_ _10886_ _10887_ VGND VGND VPWR VPWR _10888_ sky130_fd_sc_hd__xnor2_1
X_12848_ _05605_ _05606_ _05654_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__o21a_2
XFILLER_0_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15636_ _08249_ _08253_ VGND VGND VPWR VPWR _08254_ sky130_fd_sc_hd__xnor2_2
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15567_ _08176_ _08177_ VGND VGND VPWR VPWR _08188_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18355_ _10819_ _10820_ VGND VGND VPWR VPWR _10821_ sky130_fd_sc_hd__and2_1
X_12779_ _05585_ _05586_ _05563_ _05550_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__a211o_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14518_ _07198_ _07199_ _07209_ _07210_ VGND VGND VPWR VPWR _07211_ sky130_fd_sc_hd__nand4_1
X_17306_ net1050 _09266_ _09848_ _09849_ _07708_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__o221a_1
XFILLER_0_173_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15498_ _07606_ _06634_ _08136_ _07643_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18286_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[6\] _10718_ _10719_
+ VGND VGND VPWR VPWR _10753_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_86_1225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14449_ _07140_ _07141_ _07142_ VGND VGND VPWR VPWR _07144_ sky130_fd_sc_hd__a21o_1
X_17237_ _09782_ _09767_ _09769_ _05311_ VGND VGND VPWR VPWR _09784_ sky130_fd_sc_hd__o31a_1
XFILLER_0_71_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17168_ net1055 _09266_ _09716_ _09717_ _07708_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold904 top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[9\] VGND VGND
+ VPWR VPWR net1086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold915 top_inst.deskew_buff_inst.col_input\[62\] VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 top_inst.axis_out_inst.out_buff_data\[63\] VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16119_ _08700_ _08705_ _08706_ VGND VGND VPWR VPWR _08708_ sky130_fd_sc_hd__nand3_1
XFILLER_0_122_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17099_ _09647_ _09648_ _09649_ VGND VGND VPWR VPWR _09651_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19809_ _01528_ _01634_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__xor2_1
XFILLER_0_208_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22820_ _04472_ _04483_ _04484_ _04485_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22751_ top_inst.deskew_buff_inst.col_input\[122\] _05325_ VGND VGND VPWR VPWR _04422_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_211_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_91_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_220_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21702_ _03375_ _03410_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22682_ _04354_ _04355_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_1274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24421_ clknet_leaf_56_clk _00954_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21633_ _03333_ _03332_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__and2b_1
XFILLER_0_212_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24352_ clknet_leaf_24_clk _00885_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[111\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21564_ _03257_ _03259_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23303_ _04686_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__buf_2
XFILLER_0_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20515_ _02282_ _02297_ _02298_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__nand3_2
XFILLER_0_117_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24283_ clknet_leaf_10_clk _00816_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_209_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21495_ _03162_ _03187_ _03228_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23234_ _04686_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20446_ top_inst.grid_inst.data_path_wires\[16\]\[4\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[8\] VGND VGND VPWR VPWR
+ _02231_ sky130_fd_sc_hd__and3_1
XFILLER_0_244_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23165_ net78 _04687_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__or2_1
XFILLER_0_219_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20377_ _02120_ _02122_ _02162_ _02163_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_144_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22116_ _03778_ _03794_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23096_ net580 _10541_ _04646_ _04643_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22047_ _03740_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__inv_2
XFILLER_0_237_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13820_ _06526_ _06530_ _06561_ VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_214_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23998_ clknet_leaf_79_clk _00531_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_230_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13751_ _06458_ _06493_ _06421_ VGND VGND VPWR VPWR _06495_ sky130_fd_sc_hd__o21a_1
X_22949_ net413 _04557_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_82_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12702_ _05464_ _05466_ _05511_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__or3_1
X_16470_ _09007_ _09047_ VGND VGND VPWR VPWR _09048_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_1303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13682_ _06193_ _06190_ _06210_ _06208_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__and4_1
XFILLER_0_183_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15421_ _08061_ _08063_ _06734_ VGND VGND VPWR VPWR _08064_ sky130_fd_sc_hd__a21oi_1
X_12633_ _05422_ _05430_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24619_ clknet_leaf_16_clk _01152_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_127_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15352_ _07622_ _07637_ _07959_ _07958_ VGND VGND VPWR VPWR _07996_ sky130_fd_sc_hd__a31o_1
X_18140_ _10614_ _10057_ VGND VGND VPWR VPWR _10615_ sky130_fd_sc_hd__or2_1
X_12564_ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[4\] _05278_ _05282_
+ top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[3\] VGND VGND VPWR VPWR
+ _05378_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14303_ _07011_ _06996_ VGND VGND VPWR VPWR _07013_ sky130_fd_sc_hd__and2b_1
XFILLER_0_170_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18071_ _10567_ _10570_ VGND VGND VPWR VPWR _10571_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15283_ _07925_ _07928_ VGND VGND VPWR VPWR _07929_ sky130_fd_sc_hd__xor2_2
XFILLER_0_108_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12495_ _05313_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__buf_4
XFILLER_0_123_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17022_ net1118 _09575_ VGND VGND VPWR VPWR _09576_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_151_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14234_ _06825_ _06944_ VGND VGND VPWR VPWR _06946_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14165_ _06833_ _06835_ VGND VGND VPWR VPWR _06879_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13116_ top_inst.grid_inst.data_path_wires\[1\]\[4\] _05744_ _05765_ _05763_ VGND
+ VGND VPWR VPWR _05896_ sky130_fd_sc_hd__nand4_4
XFILLER_0_46_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14096_ _06809_ _06810_ VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__xnor2_2
X_18973_ _11348_ _11357_ VGND VGND VPWR VPWR _11395_ sky130_fd_sc_hd__or2b_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _05823_ _05828_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__xor2_2
X_17924_ _10377_ _10427_ VGND VGND VPWR VPWR _10429_ sky130_fd_sc_hd__or2_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17855_ _10360_ _10361_ VGND VGND VPWR VPWR _10362_ sky130_fd_sc_hd__and2_1
XFILLER_0_233_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_227_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16806_ _09193_ _09215_ _09218_ _09188_ VGND VGND VPWR VPWR _09364_ sky130_fd_sc_hd__a22o_1
XFILLER_0_234_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17786_ _10293_ VGND VGND VPWR VPWR _10294_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14998_ _07645_ _07650_ _07651_ VGND VGND VPWR VPWR _07653_ sky130_fd_sc_hd__nand3_2
X_19525_ _11688_ _11705_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__nand2_1
X_16737_ _09193_ _09188_ net217 _09210_ VGND VGND VPWR VPWR _09297_ sky130_fd_sc_hd__nand4_2
X_13949_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[2\] _06622_ _06618_
+ _06645_ VGND VGND VPWR VPWR _06669_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_53_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_73_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_241_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19456_ _01289_ _01290_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__nand2_1
X_16668_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[1\] _08183_ _09230_
+ _09231_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18407_ _10814_ _10816_ VGND VGND VPWR VPWR _10872_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15619_ _08214_ _08233_ VGND VGND VPWR VPWR _08237_ sky130_fd_sc_hd__nor2_1
X_19387_ _01195_ _01197_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__or2b_1
XFILLER_0_130_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16599_ _09159_ _09160_ _09172_ VGND VGND VPWR VPWR _09173_ sky130_fd_sc_hd__o21a_1
XFILLER_0_174_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18338_ _10579_ _10614_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[6\]
+ top_inst.grid_inst.data_path_wires\[12\]\[2\] VGND VGND VPWR VPWR _10804_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1000 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18269_ _10715_ _10735_ _10736_ VGND VGND VPWR VPWR _10737_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_1055 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20300_ _01987_ _02016_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[4\]
+ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21280_ _03006_ _03017_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold701 top_inst.deskew_buff_inst.col_input\[41\] VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold712 top_inst.deskew_buff_inst.col_input\[37\] VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold723 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[8\] VGND
+ VGND VPWR VPWR net905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20231_ _01987_ _02007_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__and3_1
XFILLER_0_188_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold734 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[9\] VGND
+ VGND VPWR VPWR net916 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold745 top_inst.axis_out_inst.out_buff_data\[80\] VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold756 top_inst.deskew_buff_inst.col_input\[71\] VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold767 top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[24\] VGND VGND
+ VPWR VPWR net949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[20\] VGND VGND
+ VPWR VPWR net960 sky130_fd_sc_hd__dlygate4sd3_1
X_20162_ _01972_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold789 top_inst.axis_in_inst.inbuf_bus\[15\] VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20093_ _01882_ _01885_ _01906_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23921_ clknet_leaf_77_clk _00454_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23852_ clknet_leaf_68_clk _00385_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_137_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22803_ _04469_ _04470_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__and2_1
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23783_ clknet_leaf_65_clk _00316_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_1227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20995_ _02761_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_64_clk clknet_4_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_16
X_22734_ _04380_ _04385_ _04404_ _06734_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22665_ _05405_ _04339_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24404_ clknet_leaf_57_clk net414 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].output_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21616_ _03346_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22596_ _04239_ _04246_ _04269_ _04223_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_69_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24335_ clknet_leaf_5_clk _00868_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_8_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21547_ _03278_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_244_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24266_ clknet_leaf_100_clk _00799_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_12280_ net756 _05164_ _05174_ _05168_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__o211a_1
XFILLER_0_244_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_209_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21478_ top_inst.grid_inst.data_path_wires\[17\]\[4\] _02897_ VGND VGND VPWR VPWR
+ _03212_ sky130_fd_sc_hd__and2b_1
XFILLER_0_181_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23217_ net102 _04714_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20429_ _02212_ _02213_ _02214_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__o21ba_1
X_24197_ clknet_leaf_15_clk _00730_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23148_ net317 _04671_ _04677_ _04675_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__o211a_1
XTAP_6211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23079_ net19 _04628_ _04637_ _04632_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__o211a_1
XTAP_5510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15970_ _08578_ _08579_ VGND VGND VPWR VPWR _08580_ sky130_fd_sc_hd__xnor2_1
XTAP_6266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsplit6 _05265_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__buf_8
XTAP_5532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14921_ net229 _07599_ _07594_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__o21a_1
XTAP_6299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold72 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[19\] VGND
+ VGND VPWR VPWR net254 sky130_fd_sc_hd__dlygate4sd3_1
X_17640_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[5\] _09496_ _10150_
+ _10151_ VGND VGND VPWR VPWR _10152_ sky130_fd_sc_hd__a22o_1
X_14852_ _07535_ _07536_ VGND VGND VPWR VPWR _07537_ sky130_fd_sc_hd__and2b_1
XTAP_5598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold83 _00158_ VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_243_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold94 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[1\]\[25\] VGND
+ VGND VPWR VPWR net276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13803_ _06507_ _06545_ VGND VGND VPWR VPWR _06546_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_230_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14783_ _07455_ _07469_ VGND VGND VPWR VPWR _07470_ sky130_fd_sc_hd__or2_1
X_17571_ _10069_ _10081_ VGND VGND VPWR VPWR _10085_ sky130_fd_sc_hd__or2b_1
XFILLER_0_187_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11995_ net760 _05004_ _05012_ _05008_ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_55_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_114_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_231_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19310_ top_inst.skew_buff_inst.row\[3\].output_reg\[7\] top_inst.axis_in_inst.inbuf_bus\[31\]
+ net34 VGND VGND VPWR VPWR _11707_ sky130_fd_sc_hd__mux2_2
XFILLER_0_86_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16522_ _09091_ _09092_ _09098_ VGND VGND VPWR VPWR _09099_ sky130_fd_sc_hd__and3_1
X_13734_ _06477_ _06478_ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19241_ _11632_ _11621_ VGND VGND VPWR VPWR _11656_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16453_ _09001_ _09002_ _09031_ VGND VGND VPWR VPWR _09032_ sky130_fd_sc_hd__o21ai_2
X_13665_ _06188_ _06214_ _06410_ VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12616_ _05385_ _05427_ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__and2_1
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15404_ _08045_ _08046_ VGND VGND VPWR VPWR _08047_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16384_ _08962_ _08963_ VGND VGND VPWR VPWR _08964_ sky130_fd_sc_hd__xnor2_1
X_19172_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[13\] _11469_ _11387_
+ VGND VGND VPWR VPWR _11589_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13596_ _06195_ _06343_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__nand2_1
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15335_ _07925_ _07928_ _07979_ VGND VGND VPWR VPWR _07980_ sky130_fd_sc_hd__a21bo_1
X_18123_ _10602_ _10057_ VGND VGND VPWR VPWR _10603_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12547_ _05357_ _05361_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_1278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_227_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15266_ _07619_ _07637_ VGND VGND VPWR VPWR _07912_ sky130_fd_sc_hd__nand2_1
X_18054_ _10525_ _10528_ _10553_ VGND VGND VPWR VPWR _10555_ sky130_fd_sc_hd__or3_1
X_12478_ _05290_ _05297_ _05299_ _05261_ VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_3 _05325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17005_ _09510_ _09512_ _09511_ VGND VGND VPWR VPWR _09559_ sky130_fd_sc_hd__a21bo_1
X_14217_ _06632_ _06650_ VGND VGND VPWR VPWR _06929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15197_ _07842_ _07844_ VGND VGND VPWR VPWR _07845_ sky130_fd_sc_hd__nor2_4
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_238_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14148_ _06856_ _06861_ VGND VGND VPWR VPWR _06862_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14079_ _06792_ _06794_ VGND VGND VPWR VPWR _06795_ sky130_fd_sc_hd__xnor2_2
X_18956_ _11375_ _11377_ _10831_ VGND VGND VPWR VPWR _11379_ sky130_fd_sc_hd__o21a_1
XFILLER_0_225_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17907_ _10296_ _10375_ _10335_ VGND VGND VPWR VPWR _10412_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_225_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18887_ _11143_ top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.weight_reg\[2\] _11309_
+ _11310_ VGND VGND VPWR VPWR _11311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_241_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17838_ _10343_ _10344_ VGND VGND VPWR VPWR _10345_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_238_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer15 _01266_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__buf_1
XFILLER_0_94_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer26 net206 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__buf_6
XFILLER_0_233_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer37 net1116 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer48 _07196_ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__buf_1
X_17769_ _10277_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_46_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_16
Xrebuffer59 _01330_ VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19508_ _01340_ _01341_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20780_ _02517_ _02548_ _02555_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19439_ _11703_ net244 _11682_ _11701_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_119_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22450_ _04103_ _04106_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21401_ top_inst.grid_inst.data_path_wires\[17\]\[4\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[5\]
+ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22381_ _04064_ _04065_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24120_ clknet_leaf_13_clk _00653_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_21332_ _03069_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_1304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24051_ clknet_leaf_34_clk _00584_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[27\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold520 top_inst.skew_buff_inst.row\[1\].has_delay.shift_reg\[0\]\[3\] VGND VGND
+ VPWR VPWR net702 sky130_fd_sc_hd__dlygate4sd3_1
X_21263_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[6\] _03000_ _03001_
+ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__and3_1
Xhold531 _00941_ VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold542 top_inst.deskew_buff_inst.col_input\[123\] VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23002_ top_inst.skew_buff_inst.row\[0\].output_reg\[2\] _04583_ VGND VGND VPWR VPWR
+ _04593_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold553 _00958_ VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__dlygate4sd3_1
X_20214_ _01993_ _11163_ _02012_ _02006_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__o211a_1
Xhold564 top_inst.skew_buff_inst.row\[3\].has_delay.shift_reg\[1\]\[5\] VGND VGND
+ VPWR VPWR net746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold575 top_inst.axis_out_inst.out_buff_data\[72\] VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__dlygate4sd3_1
X_21194_ _02923_ _02917_ _02935_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold586 top_inst.axis_out_inst.out_buff_data\[27\] VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold597 top_inst.deskew_buff_inst.col_input\[34\] VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__buf_1
XFILLER_0_198_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20145_ _01951_ _01955_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ _01871_ _01874_ _01873_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__a21o_1
XTAP_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23904_ clknet_leaf_52_clk _00437_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23835_ clknet_leaf_92_clk _00368_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clknet_4_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23766_ clknet_leaf_66_clk _00299_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_135_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11780_ net362 _04885_ _04888_ _04889_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__o211a_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20978_ _02744_ _02745_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22717_ _04092_ _04387_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23697_ clknet_leaf_121_clk net491 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13450_ _06188_ _06204_ _06209_ _06207_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__o211a_1
X_22648_ _04299_ _04302_ _04322_ _06734_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12401_ _05177_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__buf_2
X_13381_ _06152_ _06153_ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22579_ top_inst.deskew_buff_inst.col_input\[114\] _04257_ _06140_ VGND VGND VPWR
+ VPWR _04258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15120_ _07767_ _07768_ _07743_ _07744_ VGND VGND VPWR VPWR _07770_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24318_ clknet_leaf_2_clk _00851_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[93\]
+ sky130_fd_sc_hd__dfxtp_1
X_12332_ _05177_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__buf_2
XFILLER_0_105_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15051_ _07700_ _07702_ VGND VGND VPWR VPWR _07703_ sky130_fd_sc_hd__xor2_2
XFILLER_0_32_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24249_ clknet_leaf_107_clk _00782_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[40\]
+ sky130_fd_sc_hd__dfxtp_1
X_12263_ net540 _05156_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_1126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14002_ _06716_ _06719_ VGND VGND VPWR VPWR _06720_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12194_ net379 _05115_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__or2_1
Xoutput40 net40 VGND VGND VPWR VPWR output_tdata[101] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_222_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput51 net51 VGND VGND VPWR VPWR output_tdata[111] sky130_fd_sc_hd__clkbuf_4
Xoutput62 net62 VGND VGND VPWR VPWR output_tdata[121] sky130_fd_sc_hd__clkbuf_4
X_18810_ _11232_ _11235_ VGND VGND VPWR VPWR _11236_ sky130_fd_sc_hd__xor2_2
XFILLER_0_235_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput73 net73 VGND VGND VPWR VPWR output_tdata[16] sky130_fd_sc_hd__clkbuf_4
Xoutput84 net84 VGND VGND VPWR VPWR output_tdata[26] sky130_fd_sc_hd__clkbuf_4
XTAP_6041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19790_ _01599_ _01616_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput95 net95 VGND VGND VPWR VPWR output_tdata[36] sky130_fd_sc_hd__clkbuf_4
XTAP_6052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18741_ _11152_ _11132_ _11149_ _11130_ VGND VGND VPWR VPWR _11171_ sky130_fd_sc_hd__nand4_2
XTAP_6085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15953_ _08517_ _08520_ _08519_ VGND VGND VPWR VPWR _08563_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_223_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1010 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14904_ _07585_ _07586_ VGND VGND VPWR VPWR _07587_ sky130_fd_sc_hd__xnor2_1
XTAP_5373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18672_ _05787_ _11128_ _04867_ VGND VGND VPWR VPWR _11129_ sky130_fd_sc_hd__a21oi_1
XTAP_5395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ _08480_ _08481_ _08494_ VGND VGND VPWR VPWR _08496_ sky130_fd_sc_hd__nand3_1
XFILLER_0_208_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17623_ _10027_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[2\] _10115_
+ _10088_ _10052_ VGND VGND VPWR VPWR _10135_ sky130_fd_sc_hd__a32o_1
X_14835_ _07486_ _07510_ _07509_ VGND VGND VPWR VPWR _07520_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_215_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _10068_ _10069_ _06682_ VGND VGND VPWR VPWR _10070_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14766_ _07450_ _07451_ VGND VGND VPWR VPWR _07453_ sky130_fd_sc_hd__and2_1
XFILLER_0_187_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11978_ top_inst.axis_out_inst.out_buff_data\[59\] _04996_ VGND VGND VPWR VPWR _05002_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_53_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16505_ _08876_ _08677_ _09081_ VGND VGND VPWR VPWR _09082_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13717_ _06457_ _06461_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__xnor2_1
X_14697_ _07377_ _07385_ VGND VGND VPWR VPWR _07386_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_196_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17485_ _10017_ _10018_ VGND VGND VPWR VPWR _10019_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19224_ _11619_ _11638_ _11639_ _05309_ _04861_ VGND VGND VPWR VPWR _11640_ sky130_fd_sc_hd__a2111o_1
X_16436_ _09007_ _09014_ VGND VGND VPWR VPWR _09015_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13648_ _06340_ _06349_ _06394_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19155_ _11531_ _11533_ VGND VGND VPWR VPWR _11573_ sky130_fd_sc_hd__or2b_1
X_16367_ _08899_ _08902_ VGND VGND VPWR VPWR _08948_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13579_ _06297_ _06302_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18106_ _10035_ _10584_ _10590_ _10448_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__o211a_1
X_15318_ _07910_ _07912_ _07909_ VGND VGND VPWR VPWR _07963_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_82_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16298_ _08878_ _08879_ VGND VGND VPWR VPWR _08880_ sky130_fd_sc_hd__xnor2_4
X_19086_ _11427_ _11462_ _11501_ _11504_ _11500_ VGND VGND VPWR VPWR _11505_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18037_ _10521_ _10538_ VGND VGND VPWR VPWR _10539_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15249_ _07893_ _07895_ VGND VGND VPWR VPWR _07896_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1070 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19988_ _01801_ _01805_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__xor2_2
XFILLER_0_226_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18939_ _11343_ _11361_ VGND VGND VPWR VPWR _11362_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_226_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21950_ _03650_ _03646_ _03656_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20901_ _02670_ _02669_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__or2b_1
X_21881_ _03598_ _03599_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_19_clk clknet_4_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23620_ clknet_leaf_102_clk net487 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20832_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[17\] _02559_ _02578_
+ _02576_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23551_ clknet_leaf_102_clk net550 VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_20763_ _02494_ _02492_ _02510_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_193_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22502_ _05403_ _04181_ _04182_ _04183_ _05352_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__o311a_1
XFILLER_0_212_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23482_ clknet_leaf_137_clk _00015_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[72\]
+ sky130_fd_sc_hd__dfxtp_1
X_20694_ _02465_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_162_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22433_ _04058_ _04081_ _04116_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_220_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22364_ _09787_ _04047_ _04048_ _04049_ _05352_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__o311a_1
XFILLER_0_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24103_ clknet_leaf_115_clk _00636_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_143_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21315_ _03051_ _03052_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22295_ _03978_ _03981_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24034_ clknet_leaf_41_clk _00567_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold350 _01155_ VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__dlygate4sd3_1
X_21246_ _02936_ _02958_ _02985_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__o21a_1
XFILLER_0_229_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold361 _01172_ VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[6\] VGND
+ VGND VPWR VPWR net554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _00003_ VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold394 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[17\] VGND
+ VGND VPWR VPWR net576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21177_ _02907_ _02919_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_229_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_244_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20128_ _01783_ _01921_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__nor2_2
XFILLER_0_102_1176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12950_ top_inst.grid_inst.data_path_wires\[1\]\[5\] VGND VGND VPWR VPWR _05748_
+ sky130_fd_sc_hd__clkbuf_4
X_20059_ _01562_ _01872_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__nand2_1
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ net953 _04951_ _04958_ _04955_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__o211a_1
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _05685_ _05686_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__nor2_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _07308_ _07309_ _05335_ VGND VGND VPWR VPWR _07311_ sky130_fd_sc_hd__o21ai_1
X_11832_ net688 _04912_ _04919_ _04916_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__o211a_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23818_ clknet_leaf_93_clk _00351_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _07241_ _07242_ _07060_ _07064_ VGND VGND VPWR VPWR _07243_ sky130_fd_sc_hd__or4b_4
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11763_ top_inst.axis_out_inst.out_buff_data\[126\] _04877_ VGND VGND VPWR VPWR _04880_
+ sky130_fd_sc_hd__or2_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23749_ clknet_leaf_122_clk net330 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13502_ top_inst.grid_inst.data_path_wires\[2\]\[0\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[2\]\[1\]
+ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__a22o_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ _09624_ _09814_ VGND VGND VPWR VPWR _09815_ sky130_fd_sc_hd__xor2_2
X_14482_ _07083_ _07061_ _07173_ _07174_ VGND VGND VPWR VPWR _07176_ sky130_fd_sc_hd__a22oi_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16221_ _08799_ _08804_ VGND VGND VPWR VPWR _08805_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13433_ _05751_ _06192_ _06197_ _06183_ VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16152_ _08736_ _08737_ _08722_ VGND VGND VPWR VPWR _08739_ sky130_fd_sc_hd__a21o_1
XFILLER_0_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13364_ _06136_ _06137_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__nand2_1
Xrebuffer6 _09892_ VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__dlymetal6s4s_1
XFILLER_0_183_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15103_ _07747_ _07752_ VGND VGND VPWR VPWR _07753_ sky130_fd_sc_hd__xnor2_1
X_12315_ _05127_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__buf_2
X_16083_ _05755_ VGND VGND VPWR VPWR _08681_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_239_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13295_ _06068_ _06069_ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19911_ _01717_ _01732_ _07576_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__a21oi_1
X_15034_ _05887_ _07684_ _07685_ _07686_ VGND VGND VPWR VPWR _07687_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12246_ net596 _05151_ _05154_ _05155_ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19842_ _01665_ _01666_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__nor2_1
X_12177_ top_inst.axis_out_inst.out_buff_data\[16\] _05115_ VGND VGND VPWR VPWR _05116_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_102_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_208_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19773_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[13\] _01395_ _01396_
+ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16985_ _09539_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18724_ _11158_ _11150_ VGND VGND VPWR VPWR _11159_ sky130_fd_sc_hd__or2_1
XTAP_5170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15936_ _08543_ _08545_ VGND VGND VPWR VPWR _08547_ sky130_fd_sc_hd__nor2_1
XTAP_5181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_922 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18655_ _11090_ _11112_ VGND VGND VPWR VPWR _11113_ sky130_fd_sc_hd__xnor2_1
XTAP_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15867_ _08461_ _08462_ VGND VGND VPWR VPWR _08479_ sky130_fd_sc_hd__nor2_1
XTAP_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1030 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17606_ _10090_ _10097_ VGND VGND VPWR VPWR _10119_ sky130_fd_sc_hd__or2_1
XFILLER_0_235_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14818_ _07502_ _07503_ VGND VGND VPWR VPWR _07504_ sky130_fd_sc_hd__or2_1
XFILLER_0_176_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18586_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[14\] _10923_ VGND
+ VGND VPWR VPWR _11046_ sky130_fd_sc_hd__nor2_1
XTAP_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15798_ _08359_ VGND VGND VPWR VPWR _08412_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17537_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[6\] VGND VGND
+ VPWR VPWR _10056_ sky130_fd_sc_hd__buf_2
X_14749_ _07396_ _07436_ VGND VGND VPWR VPWR _07437_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17468_ _09973_ _10003_ VGND VGND VPWR VPWR _10004_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19207_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[15\] _11469_ VGND
+ VGND VPWR VPWR _11623_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16419_ _08998_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17399_ _09919_ _09917_ VGND VGND VPWR VPWR _09938_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19138_ _11551_ _11555_ VGND VGND VPWR VPWR _11556_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_144_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19069_ _11447_ _11446_ VGND VGND VPWR VPWR _11489_ sky130_fd_sc_hd__or2b_1
XFILLER_0_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_clk clknet_4_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_112_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21100_ _05317_ _02860_ _02861_ _04867_ VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__a211oi_1
X_22080_ _03770_ _03772_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_160_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21031_ _02794_ _02795_ _02784_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1042 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22982_ net992 _04575_ _04581_ _04577_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21933_ net668 _06169_ _03649_ _02909_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_1141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21864_ _03572_ _03583_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_214_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23603_ clknet_leaf_103_clk net448 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20815_ _02569_ _02571_ _02589_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__a21oi_1
X_24583_ clknet_leaf_142_clk _01116_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21795_ _03514_ _03517_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__xnor2_1
X_23534_ clknet_leaf_140_clk net669 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20746_ _02520_ _02521_ _02466_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23465_ top_inst.axis_out_inst.out_buff_data\[120\] _04864_ VGND VGND VPWR VPWR _04855_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_68_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20677_ _02389_ _02455_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22416_ top_inst.grid_inst.data_path_wires\[18\]\[7\] top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__nand2_2
XFILLER_0_66_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23396_ net62 _04658_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22347_ _04030_ _04032_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__xor2_2
XFILLER_0_104_944 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12100_ top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[1\]\[15\] _05063_
+ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13080_ _05859_ _05860_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22278_ _03897_ _03914_ _03965_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_237_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24017_ clknet_leaf_52_clk _00550_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12031_ net280 _05031_ _05032_ _05022_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold180 top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[5\] VGND
+ VGND VPWR VPWR net362 sky130_fd_sc_hd__dlygate4sd3_1
X_21229_ _02889_ _02967_ _02968_ VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__a21bo_1
Xhold191 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[9\] VGND
+ VGND VPWR VPWR net373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16770_ _09305_ _09306_ _09327_ _09328_ VGND VGND VPWR VPWR _09329_ sky130_fd_sc_hd__a211o_4
X_13982_ _05311_ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__buf_8
XFILLER_0_219_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15721_ _08289_ _08336_ VGND VGND VPWR VPWR _08337_ sky130_fd_sc_hd__nand2_1
X_12933_ _04858_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__clkbuf_8
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _10890_ _10891_ _10903_ VGND VGND VPWR VPWR _10904_ sky130_fd_sc_hd__a21oi_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _08261_ _08260_ VGND VGND VPWR VPWR _08269_ sky130_fd_sc_hd__nor2_1
X_12864_ _05616_ _05662_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14603_ _07083_ _07073_ _07291_ _07293_ VGND VGND VPWR VPWR _07294_ sky130_fd_sc_hd__nand4_1
XFILLER_0_201_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11815_ net391 _04903_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__or2_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _10827_ _10829_ _10825_ VGND VGND VPWR VPWR _10836_ sky130_fd_sc_hd__a21o_1
X_12795_ _05601_ _05602_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__xor2_1
XFILLER_0_139_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15583_ _08139_ _08157_ _08155_ _08143_ VGND VGND VPWR VPWR _08203_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17322_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[22\] _09496_ _09852_
+ _09864_ VGND VGND VPWR VPWR _09865_ sky130_fd_sc_hd__a22o_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14534_ _07226_ VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__clkbuf_1
X_11746_ _04867_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17253_ _09770_ _09776_ _09796_ _09758_ VGND VGND VPWR VPWR _09799_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14465_ net1070 _07048_ _07158_ _07159_ _06180_ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__o221a_1
XFILLER_0_126_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16204_ top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.sum_output\[5\] _08066_ _08787_
+ _08788_ VGND VGND VPWR VPWR _08789_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13416_ _05738_ _05256_ _06185_ _06183_ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17184_ _09728_ _09731_ _09732_ VGND VGND VPWR VPWR _09733_ sky130_fd_sc_hd__nand3_1
XFILLER_0_181_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14396_ _07093_ _07094_ _05336_ VGND VGND VPWR VPWR _07095_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_153_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13347_ _06084_ _06088_ _06119_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__or3_1
X_16135_ _08708_ _08719_ VGND VGND VPWR VPWR _08722_ sky130_fd_sc_hd__and2b_1
XFILLER_0_122_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16066_ top_inst.grid_inst.data_path_wires\[8\]\[3\] VGND VGND VPWR VPWR _08669_
+ sky130_fd_sc_hd__clkbuf_4
X_13278_ _06052_ _06053_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__nor2_2
XFILLER_0_110_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15017_ top_inst.grid_inst.data_path_wires\[6\]\[1\] top_inst.grid_inst.data_path_wires\[6\]\[0\]
+ _07633_ VGND VGND VPWR VPWR _07670_ sky130_fd_sc_hd__and3_1
X_12229_ net554 _05143_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__or2_1
XFILLER_0_209_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19825_ _01628_ _01626_ _01644_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19756_ _01531_ _01545_ _01544_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__a21bo_1
X_16968_ _09505_ _09521_ _09522_ VGND VGND VPWR VPWR _09523_ sky130_fd_sc_hd__and3_1
XFILLER_0_194_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18707_ top_inst.grid_inst.data_path_wires\[13\]\[7\] VGND VGND VPWR VPWR _11147_
+ sky130_fd_sc_hd__buf_4
XFILLER_0_194_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15919_ _08528_ _08529_ VGND VGND VPWR VPWR _08530_ sky130_fd_sc_hd__nand2_2
X_19687_ net253 VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__inv_2
X_16899_ _09420_ _09415_ VGND VGND VPWR VPWR _09455_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18638_ _11075_ _11073_ VGND VGND VPWR VPWR _11096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_231_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18569_ _11027_ _11029_ VGND VGND VPWR VPWR _11030_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20600_ _02351_ _02381_ _07576_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21580_ _04873_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20531_ _02275_ _02278_ net177 _02313_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_117_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23250_ net118 _04727_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20462_ _02244_ _02245_ _02193_ _02194_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_244_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22201_ _03861_ _03864_ _03862_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__a21boi_2
X_23181_ net85 _04687_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__or2_1
X_20393_ top_inst.grid_inst.data_path_wires\[16\]\[3\] top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[7\] VGND VGND VPWR VPWR
+ _02179_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22132_ _03711_ _03709_ _03682_ top_inst.grid_inst.data_path_wires\[18\]\[0\] VGND
+ VGND VPWR VPWR _03823_ sky130_fd_sc_hd__and4_1
XFILLER_0_219_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1030 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22063_ _03311_ _03756_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__and2_1
XTAP_6629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21014_ top_inst.deskew_buff_inst.col_input\[58\] _11723_ _02763_ _02780_ VGND VGND
+ VPWR VPWR _02781_ sky130_fd_sc_hd__a22o_1
XFILLER_0_227_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22965_ top_inst.skew_buff_inst.row\[1\].output_reg\[2\] _04570_ VGND VGND VPWR VPWR
+ _04572_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21916_ _03631_ _03632_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22896_ net784 _04522_ _04532_ _04524_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24635_ clknet_leaf_24_clk _01168_ VGND VGND VPWR VPWR top_inst.axis_out_inst.out_buff_data\[111\]
+ sky130_fd_sc_hd__dfxtp_1
X_21847_ _03566_ _03567_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__and2_1
XFILLER_0_183_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12580_ _05391_ _05393_ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__xnor2_1
X_24566_ clknet_leaf_137_clk _01099_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_148_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21778_ _03472_ _03479_ _03497_ _03452_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_38_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23517_ clknet_leaf_138_clk net754 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[2\].delayed_pass.shift_reg\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_20729_ _02459_ _02481_ _02480_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24497_ clknet_leaf_108_clk _01030_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_110_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14250_ _06931_ _06930_ VGND VGND VPWR VPWR _06961_ sky130_fd_sc_hd__or2b_1
XFILLER_0_123_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23448_ net654 _04840_ _04846_ _04844_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13201_ _05977_ _05978_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__nor2_1
X_14181_ _06650_ _06630_ VGND VGND VPWR VPWR _06894_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23379_ net710 _04804_ _04809_ _04808_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13132_ _05853_ _05862_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_237_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13063_ _05818_ _05843_ _05399_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17940_ _10443_ _10444_ VGND VGND VPWR VPWR _10445_ sky130_fd_sc_hd__and2_1
X_12014_ _05009_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__clkbuf_2
X_17871_ _10296_ _10376_ VGND VGND VPWR VPWR _10377_ sky130_fd_sc_hd__xnor2_4
X_19610_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[3\] _11704_ _11708_
+ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16822_ _09376_ _09378_ _09379_ VGND VGND VPWR VPWR _09380_ sky130_fd_sc_hd__nand3_1
XFILLER_0_219_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19541_ _01371_ _01372_ _01373_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__nand3_2
X_16753_ _09282_ _09311_ _09312_ VGND VGND VPWR VPWR _09313_ sky130_fd_sc_hd__nor3_2
XFILLER_0_219_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13965_ net1072 _06660_ _06683_ _06684_ VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__o211a_1
XFILLER_0_232_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15704_ _08147_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.weight_reg\[2\] _08317_
+ _08318_ VGND VGND VPWR VPWR _08320_ sky130_fd_sc_hd__nand4_2
X_12916_ _05699_ _05720_ _05440_ VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_198_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19472_ _01299_ _01305_ VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__xnor2_1
X_16684_ _09246_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_216_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13896_ top_inst.grid_inst.data_path_wires\[3\]\[5\] VGND VGND VPWR VPWR _06630_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18423_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[10\] _10793_ VGND
+ VGND VPWR VPWR _10887_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15635_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[5\] _08252_ VGND
+ VGND VPWR VPWR _08253_ sky130_fd_sc_hd__xor2_2
X_12847_ _05280_ _05273_ _05306_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18354_ _10776_ _10751_ VGND VGND VPWR VPWR _10820_ sky130_fd_sc_hd__or2b_1
XFILLER_0_186_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15566_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[2\] _08186_ VGND
+ VGND VPWR VPWR _08187_ sky130_fd_sc_hd__xor2_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12778_ _05563_ _05550_ _05585_ _05586_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_17_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17305_ _09830_ _09831_ _09847_ _07439_ VGND VGND VPWR VPWR _09849_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14517_ _07207_ _07208_ _07175_ VGND VGND VPWR VPWR _07210_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18285_ _10724_ _10733_ _10735_ VGND VGND VPWR VPWR _10752_ sky130_fd_sc_hd__o21ai_1
X_15497_ _08135_ _06620_ VGND VGND VPWR VPWR _08136_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17236_ _09767_ _09769_ _09782_ VGND VGND VPWR VPWR _09783_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_153_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14448_ _07140_ _07141_ _07142_ VGND VGND VPWR VPWR _07143_ sky130_fd_sc_hd__nand3_1
XFILLER_0_43_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17167_ _09697_ _09715_ _06178_ VGND VGND VPWR VPWR _09717_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14379_ top_inst.skew_buff_inst.row\[1\].output_reg\[5\] top_inst.axis_in_inst.inbuf_bus\[13\]
+ net208 VGND VGND VPWR VPWR _07081_ sky130_fd_sc_hd__mux2_4
Xhold905 top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.sum_output\[2\] VGND VGND
+ VPWR VPWR net1087 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold916 top_inst.deskew_buff_inst.col_input\[27\] VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold927 top_inst.axis_in_inst.inbuf_bus\[21\] VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16118_ _08705_ _08706_ _08700_ VGND VGND VPWR VPWR _08707_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17098_ _09647_ _09648_ _09649_ VGND VGND VPWR VPWR _09650_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16049_ _08652_ _08655_ VGND VGND VPWR VPWR _08656_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_177_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19808_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[15\] _01480_ VGND
+ VGND VPWR VPWR _01634_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19739_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[13\] _01480_ VGND
+ VGND VPWR VPWR _01567_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_233_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22750_ _04401_ _04419_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__nand2_2
XFILLER_0_95_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21701_ _03423_ _03427_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_177_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22681_ _04352_ _04353_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24420_ clknet_leaf_58_clk _00953_ VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21632_ _03348_ _03361_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_133_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24351_ clknet_leaf_26_clk _00884_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[110\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21563_ _03210_ _03294_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_168_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23302_ _04684_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_191_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20514_ _02294_ _02295_ _02296_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24282_ clknet_leaf_13_clk _00815_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_244_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21494_ _03184_ _03186_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__nor2_1
XFILLER_0_244_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23233_ _04684_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20445_ top_inst.grid_inst.data_path_wires\[16\]\[4\] _02015_ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[8\]
+ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_160_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23164_ _04686_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__buf_2
X_20376_ _02160_ _02161_ _02143_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22115_ _03799_ _03798_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__nor2_1
XTAP_6404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23095_ net624 _05323_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__or2_1
XTAP_6426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22046_ _03705_ _03703_ _03682_ _03680_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__and4_2
XTAP_6459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23997_ clknet_leaf_79_clk _00530_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[3\].pe_inst.weight_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13750_ _06421_ _06458_ _06493_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__nor3_1
X_22948_ _10583_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__clkbuf_4
X_12701_ _05464_ _05466_ _05511_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_74_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13681_ _06423_ _06426_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__xnor2_1
X_22879_ net746 _04517_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_1364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15420_ _08022_ _08024_ _08062_ VGND VGND VPWR VPWR _08063_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_13_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12632_ _05412_ _05421_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24618_ clknet_leaf_21_clk _01151_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_38_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12563_ _05298_ _05272_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__nand2_1
X_15351_ _07990_ _07994_ VGND VGND VPWR VPWR _07995_ sky130_fd_sc_hd__xor2_1
XFILLER_0_38_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24549_ clknet_leaf_131_clk _01082_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_54_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14302_ _06996_ _07011_ VGND VGND VPWR VPWR _07012_ sky130_fd_sc_hd__and2b_1
XFILLER_0_227_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18070_ _10568_ _10569_ VGND VGND VPWR VPWR _10570_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15282_ _07926_ _07927_ VGND VGND VPWR VPWR _07928_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12494_ _05312_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__buf_12
XFILLER_0_81_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17021_ _09573_ _09574_ VGND VGND VPWR VPWR _09575_ sky130_fd_sc_hd__xnor2_2
X_14233_ _06825_ _06944_ VGND VGND VPWR VPWR _06945_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14164_ _06875_ _06877_ VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13115_ _05744_ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[3\]
+ top_inst.grid_inst.data_path_wires\[1\]\[4\] VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14095_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.weight_reg\[5\] _06626_ VGND
+ VGND VPWR VPWR _06810_ sky130_fd_sc_hd__nand2_1
X_18972_ _11356_ _11354_ VGND VGND VPWR VPWR _11394_ sky130_fd_sc_hd__or2b_1
XFILLER_0_237_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13046_ _05826_ _05827_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__xor2_2
X_17923_ _10377_ _10427_ VGND VGND VPWR VPWR _10428_ sky130_fd_sc_hd__nand2_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17854_ _10324_ _10359_ VGND VGND VPWR VPWR _10361_ sky130_fd_sc_hd__or2_1
XFILLER_0_205_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16805_ _09334_ _09335_ VGND VGND VPWR VPWR _09363_ sky130_fd_sc_hd__nand2_1
X_17785_ top_inst.grid_inst.data_path_wires\[11\]\[6\] top_inst.grid_inst.data_path_wires\[11\]\[5\]
+ top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[4\] top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.weight_reg\[3\]
+ VGND VGND VPWR VPWR _10293_ sky130_fd_sc_hd__and4_1
XFILLER_0_227_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14997_ _07650_ _07651_ _07645_ VGND VGND VPWR VPWR _07652_ sky130_fd_sc_hd__a21o_1
XFILLER_0_221_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19524_ _01350_ _01356_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__xor2_1
XFILLER_0_233_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16736_ _09193_ net216 _09209_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _09296_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13948_ top_inst.grid_inst.rows\[0\].cols\[3\].pe_inst.sum_output\[2\] _06660_ _06668_
+ _06639_ VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19455_ _01221_ _01259_ _01287_ _01288_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__o22ai_2
X_16667_ _07617_ VGND VGND VPWR VPWR _09231_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13879_ top_inst.grid_inst.data_path_wires\[3\]\[0\] VGND VGND VPWR VPWR _06618_
+ sky130_fd_sc_hd__buf_2
XFILLER_0_201_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18406_ _10839_ _10870_ VGND VGND VPWR VPWR _10871_ sky130_fd_sc_hd__xor2_1
XFILLER_0_243_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15618_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[4\] _07048_ _08235_
+ _08236_ _07708_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__o221a_1
X_19386_ _01221_ _01222_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16598_ _09150_ _09158_ VGND VGND VPWR VPWR _09172_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18337_ top_inst.grid_inst.data_path_wires\[12\]\[2\] _10579_ _10614_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[6\]
+ VGND VGND VPWR VPWR _10803_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15549_ _08135_ _08155_ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[0\]
+ VGND VGND VPWR VPWR _08172_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18268_ _10723_ _10734_ VGND VGND VPWR VPWR _10736_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_942 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17219_ net1022 _09266_ _09765_ _09766_ _07708_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__o221a_1
XFILLER_0_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1067 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18199_ top_inst.grid_inst.rows\[1\].cols\[2\].pe_inst.sum_output\[3\] _10648_ _10649_
+ VGND VGND VPWR VPWR _10669_ sky130_fd_sc_hd__a21bo_1
Xhold702 top_inst.deskew_buff_inst.col_input\[118\] VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[27\] VGND
+ VGND VPWR VPWR net895 sky130_fd_sc_hd__dlygate4sd3_1
X_20230_ _02004_ _11163_ _02023_ _02006_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold724 top_inst.deskew_buff_inst.col_input\[26\] VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__buf_1
Xhold735 top_inst.deskew_buff_inst.col_input\[0\] VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[19\] VGND VGND
+ VPWR VPWR net928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold757 top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.sum_output\[19\] VGND VGND
+ VPWR VPWR net939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[0\] VGND VGND
+ VPWR VPWR net950 sky130_fd_sc_hd__dlygate4sd3_1
X_20161_ _11722_ _01971_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__and2_4
XFILLER_0_12_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold779 top_inst.grid_inst.rows\[2\].cols\[1\].pe_inst.sum_output\[21\] VGND VGND
+ VPWR VPWR net961 sky130_fd_sc_hd__dlygate4sd3_1
X_20092_ _01879_ _01905_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_244_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23920_ clknet_leaf_76_clk _00453_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_97_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23851_ clknet_leaf_68_clk _00384_ VGND VGND VPWR VPWR top_inst.grid_inst.data_path_wires\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_237_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22802_ _04388_ _04446_ _04468_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__nand3_1
XFILLER_0_170_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23782_ clknet_leaf_65_clk _00315_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.sum_output\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20994_ _02730_ _02733_ _02756_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__a21oi_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22733_ _04380_ _04385_ _04404_ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_211_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22664_ _04337_ _04338_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24403_ clknet_leaf_55_clk net767 VGND VGND VPWR VPWR top_inst.skew_buff_inst.row\[2\].output_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21615_ _03311_ _03345_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__and2_1
X_22595_ _04271_ _04272_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21546_ _03246_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__buf_2
X_24334_ clknet_leaf_5_clk _00867_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[3\].cols\[3\].pe_inst.weight_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_117_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_836 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24265_ clknet_leaf_101_clk _00798_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21477_ top_inst.grid_inst.data_path_wires\[17\]\[6\] top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[5\]
+ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__nand2_1
XFILLER_0_205_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23216_ net822 _04713_ _04716_ _04717_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20428_ _02125_ _02168_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__nor2_1
X_24196_ clknet_leaf_15_clk _00729_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1010 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23147_ net70 _04672_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20359_ top_inst.grid_inst.data_path_wires\[16\]\[6\] _01986_ _02020_ top_inst.grid_inst.rows\[3\].cols\[1\].pe_inst.weight_reg\[0\]
+ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__and4_1
XTAP_6201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23078_ top_inst.axis_in_inst.inbuf_bus\[26\] _04629_ VGND VGND VPWR VPWR _04637_
+ sky130_fd_sc_hd__or2_1
XTAP_5500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14920_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[20\] _07595_ VGND
+ VGND VPWR VPWR _07599_ sky130_fd_sc_hd__and2_1
XTAP_5533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22029_ net581 _06169_ _03724_ _03702_ VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__o211a_1
XTAP_6289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14851_ _07527_ _07502_ _07534_ VGND VGND VPWR VPWR _07536_ sky130_fd_sc_hd__or3b_1
XTAP_5588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold73 _00154_ VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold84 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[28\] VGND
+ VGND VPWR VPWR net266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_230_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold95 _00288_ VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13802_ _06543_ _06544_ VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_216_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17570_ _10071_ _10082_ _10084_ _10049_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__o211a_1
X_14782_ _07467_ _07468_ VGND VGND VPWR VPWR _07469_ sky130_fd_sc_hd__nand2_1
XTAP_4898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11994_ net447 _05010_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__or2_1
XFILLER_0_187_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16521_ _09093_ _09097_ VGND VGND VPWR VPWR _09098_ sky130_fd_sc_hd__xor2_1
XFILLER_0_168_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13733_ _06474_ _06476_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_230_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19240_ _11653_ _11654_ VGND VGND VPWR VPWR _11655_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16452_ _09028_ _09030_ VGND VGND VPWR VPWR _09031_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13664_ top_inst.grid_inst.data_path_wires\[2\]\[2\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[7\]
+ VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15403_ _08005_ _08044_ VGND VGND VPWR VPWR _08046_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12615_ _05385_ _05427_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__nor2_1
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19171_ _11556_ _11571_ _11569_ VGND VGND VPWR VPWR _11588_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16383_ _08695_ _08673_ VGND VGND VPWR VPWR _08963_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13595_ top_inst.grid_inst.data_path_wires\[2\]\[7\] top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[1\]
+ top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.weight_reg\[0\] VGND VGND VPWR VPWR
+ _06343_ sky130_fd_sc_hd__and3_1
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18122_ top_inst.grid_inst.rows\[2\].cols\[2\].pe_inst.weight_reg\[2\] VGND VGND
+ VPWR VPWR _10602_ sky130_fd_sc_hd__buf_4
XFILLER_0_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15334_ _07927_ _07926_ VGND VGND VPWR VPWR _07979_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12546_ _05339_ _05360_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18053_ _10525_ _10528_ _10553_ VGND VGND VPWR VPWR _10554_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15265_ _07909_ _07910_ VGND VGND VPWR VPWR _07911_ sky130_fd_sc_hd__nor2_1
X_12477_ _05298_ _05294_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__or2_1
X_17004_ _09555_ _09556_ _09554_ VGND VGND VPWR VPWR _09558_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 _06178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_227_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14216_ _06926_ _06927_ VGND VGND VPWR VPWR _06928_ sky130_fd_sc_hd__nor2_1
X_15196_ _07843_ VGND VGND VPWR VPWR _07844_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14147_ _06859_ _06860_ VGND VGND VPWR VPWR _06861_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14078_ _06749_ _06755_ _06793_ VGND VGND VPWR VPWR _06794_ sky130_fd_sc_hd__o21ai_2
X_18955_ _11375_ _11377_ VGND VGND VPWR VPWR _11378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_238_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13029_ top_inst.grid_inst.data_path_wires\[1\]\[0\] top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[4\]
+ top_inst.grid_inst.rows\[0\].cols\[1\].pe_inst.weight_reg\[3\] top_inst.grid_inst.data_path_wires\[1\]\[1\]
+ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__a22o_1
X_17906_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[11\] _10367_ _10283_
+ VGND VGND VPWR VPWR _10411_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18886_ _11158_ top_inst.grid_inst.data_path_wires\[13\]\[4\] _11156_ _11138_ VGND
+ VGND VPWR VPWR _11310_ sky130_fd_sc_hd__nand4_2
XFILLER_0_158_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17837_ _10298_ _10301_ _10299_ VGND VGND VPWR VPWR _10344_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_59_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_240_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer16 net197 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_1
Xrebuffer27 _07167_ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer38 _09514_ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_1
X_17768_ _09661_ _10276_ VGND VGND VPWR VPWR _10277_ sky130_fd_sc_hd__and2_1
Xrebuffer49 _01262_ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16719_ _09273_ _09278_ _09279_ VGND VGND VPWR VPWR _09280_ sky130_fd_sc_hd__nand3_2
XFILLER_0_159_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19507_ _01290_ _01293_ _01289_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_92_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17699_ _10207_ _10208_ VGND VGND VPWR VPWR _10209_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19438_ top_inst.grid_inst.rows\[3\].cols\[0\].pe_inst.weight_reg\[2\] _11696_ _01270_
+ _01271_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_1212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19369_ _01203_ _01204_ top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[4\]
+ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21400_ _03134_ _03135_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22380_ _04059_ _04063_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21331_ _02135_ _03068_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24050_ clknet_leaf_34_clk _00583_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[0\].pe_inst.sum_output\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold510 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[2\]\[14\] VGND
+ VGND VPWR VPWR net692 sky130_fd_sc_hd__dlygate4sd3_1
X_21262_ top_inst.grid_inst.data_path_wires\[17\]\[6\] top_inst.grid_inst.data_path_wires\[17\]\[5\]
+ top_inst.grid_inst.rows\[3\].cols\[2\].pe_inst.weight_reg\[1\] _02882_ VGND VGND
+ VPWR VPWR _03001_ sky130_fd_sc_hd__nand4_1
XFILLER_0_13_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold521 _00961_ VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23001_ net983 _04588_ _04592_ _04590_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__o211a_1
Xhold532 top_inst.axis_out_inst.out_buff_data\[109\] VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold543 top_inst.axis_out_inst.out_buff_data\[114\] VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__dlygate4sd3_1
X_20213_ _02011_ _11689_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__or2_1
Xhold554 top_inst.axis_out_inst.out_buff_data\[29\] VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold565 top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[26\] VGND
+ VGND VPWR VPWR net747 sky130_fd_sc_hd__dlygate4sd3_1
X_21193_ _02927_ _02934_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_198_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold576 top_inst.deskew_buff_inst.col_input\[35\] VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold587 top_inst.skew_buff_inst.row\[2\].has_delay.shift_reg\[1\]\[1\] VGND VGND
+ VPWR VPWR net769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20144_ _01953_ _01954_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__nor2_1
Xhold598 top_inst.deskew_buff_inst.row\[1\].delayed_pass.shift_reg\[0\]\[4\] VGND
+ VGND VPWR VPWR net780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20075_ _01889_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__clkbuf_1
XTAP_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23903_ clknet_leaf_59_clk _00436_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23834_ clknet_leaf_92_clk _00367_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[2\].pe_inst.sum_output\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23765_ clknet_leaf_66_clk _00298_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[0\].cols\[0\].pe_inst.weight_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_20977_ _02742_ _02743_ _02473_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_212_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22716_ _04218_ _04387_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__or2_2
XFILLER_0_113_1432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23696_ clknet_leaf_120_clk net401 VGND VGND VPWR VPWR top_inst.deskew_buff_inst.row\[0\].delayed_pass.shift_reg\[0\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22647_ _04299_ _04302_ _04322_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12400_ net480 _05230_ _05242_ _05234_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__o211a_1
X_13380_ _06120_ _06123_ _06151_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__and3_1
X_22578_ _04253_ _04256_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24317_ clknet_leaf_1_clk _00850_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[92\]
+ sky130_fd_sc_hd__dfxtp_1
X_12331_ net811 _05191_ _05203_ _05195_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21529_ _03215_ _03217_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__and2_1
XFILLER_0_181_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15050_ _07677_ _07678_ _07701_ VGND VGND VPWR VPWR _07702_ sky130_fd_sc_hd__o21ai_2
X_12262_ _05044_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__buf_2
XFILLER_0_133_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24248_ clknet_leaf_108_clk _00781_ VGND VGND VPWR VPWR top_inst.deskew_buff_inst.col_input\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14001_ _06717_ _06718_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24179_ clknet_leaf_29_clk _00712_ VGND VGND VPWR VPWR top_inst.grid_inst.rows\[2\].cols\[3\].pe_inst.sum_output\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12193_ net365 _05123_ _05124_ _05114_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput41 net41 VGND VGND VPWR VPWR output_tdata[102] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput52 net52 VGND VGND VPWR VPWR output_tdata[112] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_1403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput63 net63 VGND VGND VPWR VPWR output_tdata[122] sky130_fd_sc_hd__clkbuf_4
Xoutput74 net74 VGND VGND VPWR VPWR output_tdata[17] sky130_fd_sc_hd__clkbuf_4
XTAP_6031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput85 net85 VGND VGND VPWR VPWR output_tdata[27] sky130_fd_sc_hd__clkbuf_4
XTAP_6053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput96 net96 VGND VGND VPWR VPWR output_tdata[37] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18740_ _11132_ _11149_ _11130_ _11152_ VGND VGND VPWR VPWR _11170_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15952_ _08517_ _08561_ VGND VGND VPWR VPWR _08562_ sky130_fd_sc_hd__xnor2_1
XTAP_6075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14903_ _07531_ _07530_ _07564_ _07582_ VGND VGND VPWR VPWR _07586_ sky130_fd_sc_hd__o2bb2a_1
XTAP_5363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18671_ _11097_ _11113_ _11126_ _11127_ VGND VGND VPWR VPWR _11128_ sky130_fd_sc_hd__a211o_1
XFILLER_0_222_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ _08480_ _08481_ _08494_ VGND VGND VPWR VPWR _08495_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_203_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_215_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17622_ top_inst.grid_inst.rows\[1\].cols\[1\].pe_inst.sum_output\[4\] _10107_ _10108_
+ VGND VGND VPWR VPWR _10134_ sky130_fd_sc_hd__a21boi_2
X_14834_ net1066 _07048_ _07518_ _07519_ _06180_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__o221a_1
XTAP_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17553_ _10061_ _10066_ _10067_ VGND VGND VPWR VPWR _10069_ sky130_fd_sc_hd__nand3_2
X_14765_ _07450_ _07451_ VGND VGND VPWR VPWR _07452_ sky130_fd_sc_hd__nor2_1
XTAP_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ net973 _04990_ _05001_ _04995_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16504_ _08679_ _08697_ VGND VGND VPWR VPWR _09081_ sky130_fd_sc_hd__nand2_1
X_13716_ _06421_ _06460_ VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__xnor2_1
X_17484_ top_inst.grid_inst.rows\[1\].cols\[0\].pe_inst.sum_output\[31\] _10005_ VGND
+ VGND VPWR VPWR _10018_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14696_ _07383_ _07384_ VGND VGND VPWR VPWR _07385_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19223_ _11619_ _11638_ VGND VGND VPWR VPWR _11639_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16435_ _09012_ _09013_ VGND VGND VPWR VPWR _09014_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13647_ _06327_ _06339_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19154_ _11556_ _11571_ VGND VGND VPWR VPWR _11572_ sky130_fd_sc_hd__xor2_2
XFILLER_0_26_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16366_ _08944_ _08946_ VGND VGND VPWR VPWR _08947_ sky130_fd_sc_hd__xnor2_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13578_ _06326_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18105_ _10589_ _08674_ VGND VGND VPWR VPWR _10590_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15317_ _07960_ _07961_ VGND VGND VPWR VPWR _07962_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_895 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12529_ _05340_ _05344_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19085_ _11457_ _11460_ VGND VGND VPWR VPWR _11504_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16297_ _08695_ _08669_ VGND VGND VPWR VPWR _08879_ sky130_fd_sc_hd__nand2_2
XFILLER_0_124_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18036_ _10536_ _10537_ VGND VGND VPWR VPWR _10538_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15248_ _07840_ _07852_ _07894_ VGND VGND VPWR VPWR _07895_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15179_ _07613_ _07637_ VGND VGND VPWR VPWR _07827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_239_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19987_ _01803_ _01804_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__and2b_1
XFILLER_0_123_1082 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18938_ _11358_ _11360_ VGND VGND VPWR VPWR _11361_ sky130_fd_sc_hd__xnor2_1
.ends

