module top_hardened (clk,
    input_tready,
    input_tvalid,
    load_weight,
    output_tready,
    output_tvalid,
    reset,
    input_tdata,
    output_tdata);
 input clk;
 output input_tready;
 input input_tvalid;
 input load_weight;
 input output_tready;
 output output_tvalid;
 input reset;
 input [31:0] input_tdata;
 output [127:0] output_tdata;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire \top_inst.axis_in_inst.inbuf_bus[0] ;
 wire \top_inst.axis_in_inst.inbuf_bus[10] ;
 wire \top_inst.axis_in_inst.inbuf_bus[11] ;
 wire \top_inst.axis_in_inst.inbuf_bus[12] ;
 wire \top_inst.axis_in_inst.inbuf_bus[13] ;
 wire \top_inst.axis_in_inst.inbuf_bus[14] ;
 wire \top_inst.axis_in_inst.inbuf_bus[15] ;
 wire \top_inst.axis_in_inst.inbuf_bus[16] ;
 wire \top_inst.axis_in_inst.inbuf_bus[17] ;
 wire \top_inst.axis_in_inst.inbuf_bus[18] ;
 wire \top_inst.axis_in_inst.inbuf_bus[19] ;
 wire \top_inst.axis_in_inst.inbuf_bus[1] ;
 wire \top_inst.axis_in_inst.inbuf_bus[20] ;
 wire \top_inst.axis_in_inst.inbuf_bus[21] ;
 wire \top_inst.axis_in_inst.inbuf_bus[22] ;
 wire \top_inst.axis_in_inst.inbuf_bus[23] ;
 wire \top_inst.axis_in_inst.inbuf_bus[24] ;
 wire \top_inst.axis_in_inst.inbuf_bus[25] ;
 wire \top_inst.axis_in_inst.inbuf_bus[26] ;
 wire \top_inst.axis_in_inst.inbuf_bus[27] ;
 wire \top_inst.axis_in_inst.inbuf_bus[28] ;
 wire \top_inst.axis_in_inst.inbuf_bus[29] ;
 wire \top_inst.axis_in_inst.inbuf_bus[2] ;
 wire \top_inst.axis_in_inst.inbuf_bus[30] ;
 wire \top_inst.axis_in_inst.inbuf_bus[31] ;
 wire \top_inst.axis_in_inst.inbuf_bus[3] ;
 wire \top_inst.axis_in_inst.inbuf_bus[4] ;
 wire \top_inst.axis_in_inst.inbuf_bus[5] ;
 wire \top_inst.axis_in_inst.inbuf_bus[6] ;
 wire \top_inst.axis_in_inst.inbuf_bus[7] ;
 wire \top_inst.axis_in_inst.inbuf_bus[8] ;
 wire \top_inst.axis_in_inst.inbuf_bus[9] ;
 wire \top_inst.axis_in_inst.inbuf_valid ;
 wire \top_inst.axis_out_inst.out_buff_data[0] ;
 wire \top_inst.axis_out_inst.out_buff_data[100] ;
 wire \top_inst.axis_out_inst.out_buff_data[101] ;
 wire \top_inst.axis_out_inst.out_buff_data[102] ;
 wire \top_inst.axis_out_inst.out_buff_data[103] ;
 wire \top_inst.axis_out_inst.out_buff_data[104] ;
 wire \top_inst.axis_out_inst.out_buff_data[105] ;
 wire \top_inst.axis_out_inst.out_buff_data[106] ;
 wire \top_inst.axis_out_inst.out_buff_data[107] ;
 wire \top_inst.axis_out_inst.out_buff_data[108] ;
 wire \top_inst.axis_out_inst.out_buff_data[109] ;
 wire \top_inst.axis_out_inst.out_buff_data[10] ;
 wire \top_inst.axis_out_inst.out_buff_data[110] ;
 wire \top_inst.axis_out_inst.out_buff_data[111] ;
 wire \top_inst.axis_out_inst.out_buff_data[112] ;
 wire \top_inst.axis_out_inst.out_buff_data[113] ;
 wire \top_inst.axis_out_inst.out_buff_data[114] ;
 wire \top_inst.axis_out_inst.out_buff_data[115] ;
 wire \top_inst.axis_out_inst.out_buff_data[116] ;
 wire \top_inst.axis_out_inst.out_buff_data[117] ;
 wire \top_inst.axis_out_inst.out_buff_data[118] ;
 wire \top_inst.axis_out_inst.out_buff_data[119] ;
 wire \top_inst.axis_out_inst.out_buff_data[11] ;
 wire \top_inst.axis_out_inst.out_buff_data[120] ;
 wire \top_inst.axis_out_inst.out_buff_data[121] ;
 wire \top_inst.axis_out_inst.out_buff_data[122] ;
 wire \top_inst.axis_out_inst.out_buff_data[123] ;
 wire \top_inst.axis_out_inst.out_buff_data[124] ;
 wire \top_inst.axis_out_inst.out_buff_data[125] ;
 wire \top_inst.axis_out_inst.out_buff_data[126] ;
 wire \top_inst.axis_out_inst.out_buff_data[127] ;
 wire \top_inst.axis_out_inst.out_buff_data[12] ;
 wire \top_inst.axis_out_inst.out_buff_data[13] ;
 wire \top_inst.axis_out_inst.out_buff_data[14] ;
 wire \top_inst.axis_out_inst.out_buff_data[15] ;
 wire \top_inst.axis_out_inst.out_buff_data[16] ;
 wire \top_inst.axis_out_inst.out_buff_data[17] ;
 wire \top_inst.axis_out_inst.out_buff_data[18] ;
 wire \top_inst.axis_out_inst.out_buff_data[19] ;
 wire \top_inst.axis_out_inst.out_buff_data[1] ;
 wire \top_inst.axis_out_inst.out_buff_data[20] ;
 wire \top_inst.axis_out_inst.out_buff_data[21] ;
 wire \top_inst.axis_out_inst.out_buff_data[22] ;
 wire \top_inst.axis_out_inst.out_buff_data[23] ;
 wire \top_inst.axis_out_inst.out_buff_data[24] ;
 wire \top_inst.axis_out_inst.out_buff_data[25] ;
 wire \top_inst.axis_out_inst.out_buff_data[26] ;
 wire \top_inst.axis_out_inst.out_buff_data[27] ;
 wire \top_inst.axis_out_inst.out_buff_data[28] ;
 wire \top_inst.axis_out_inst.out_buff_data[29] ;
 wire \top_inst.axis_out_inst.out_buff_data[2] ;
 wire \top_inst.axis_out_inst.out_buff_data[30] ;
 wire \top_inst.axis_out_inst.out_buff_data[31] ;
 wire \top_inst.axis_out_inst.out_buff_data[32] ;
 wire \top_inst.axis_out_inst.out_buff_data[33] ;
 wire \top_inst.axis_out_inst.out_buff_data[34] ;
 wire \top_inst.axis_out_inst.out_buff_data[35] ;
 wire \top_inst.axis_out_inst.out_buff_data[36] ;
 wire \top_inst.axis_out_inst.out_buff_data[37] ;
 wire \top_inst.axis_out_inst.out_buff_data[38] ;
 wire \top_inst.axis_out_inst.out_buff_data[39] ;
 wire \top_inst.axis_out_inst.out_buff_data[3] ;
 wire \top_inst.axis_out_inst.out_buff_data[40] ;
 wire \top_inst.axis_out_inst.out_buff_data[41] ;
 wire \top_inst.axis_out_inst.out_buff_data[42] ;
 wire \top_inst.axis_out_inst.out_buff_data[43] ;
 wire \top_inst.axis_out_inst.out_buff_data[44] ;
 wire \top_inst.axis_out_inst.out_buff_data[45] ;
 wire \top_inst.axis_out_inst.out_buff_data[46] ;
 wire \top_inst.axis_out_inst.out_buff_data[47] ;
 wire \top_inst.axis_out_inst.out_buff_data[48] ;
 wire \top_inst.axis_out_inst.out_buff_data[49] ;
 wire \top_inst.axis_out_inst.out_buff_data[4] ;
 wire \top_inst.axis_out_inst.out_buff_data[50] ;
 wire \top_inst.axis_out_inst.out_buff_data[51] ;
 wire \top_inst.axis_out_inst.out_buff_data[52] ;
 wire \top_inst.axis_out_inst.out_buff_data[53] ;
 wire \top_inst.axis_out_inst.out_buff_data[54] ;
 wire \top_inst.axis_out_inst.out_buff_data[55] ;
 wire \top_inst.axis_out_inst.out_buff_data[56] ;
 wire \top_inst.axis_out_inst.out_buff_data[57] ;
 wire \top_inst.axis_out_inst.out_buff_data[58] ;
 wire \top_inst.axis_out_inst.out_buff_data[59] ;
 wire \top_inst.axis_out_inst.out_buff_data[5] ;
 wire \top_inst.axis_out_inst.out_buff_data[60] ;
 wire \top_inst.axis_out_inst.out_buff_data[61] ;
 wire \top_inst.axis_out_inst.out_buff_data[62] ;
 wire \top_inst.axis_out_inst.out_buff_data[63] ;
 wire \top_inst.axis_out_inst.out_buff_data[64] ;
 wire \top_inst.axis_out_inst.out_buff_data[65] ;
 wire \top_inst.axis_out_inst.out_buff_data[66] ;
 wire \top_inst.axis_out_inst.out_buff_data[67] ;
 wire \top_inst.axis_out_inst.out_buff_data[68] ;
 wire \top_inst.axis_out_inst.out_buff_data[69] ;
 wire \top_inst.axis_out_inst.out_buff_data[6] ;
 wire \top_inst.axis_out_inst.out_buff_data[70] ;
 wire \top_inst.axis_out_inst.out_buff_data[71] ;
 wire \top_inst.axis_out_inst.out_buff_data[72] ;
 wire \top_inst.axis_out_inst.out_buff_data[73] ;
 wire \top_inst.axis_out_inst.out_buff_data[74] ;
 wire \top_inst.axis_out_inst.out_buff_data[75] ;
 wire \top_inst.axis_out_inst.out_buff_data[76] ;
 wire \top_inst.axis_out_inst.out_buff_data[77] ;
 wire \top_inst.axis_out_inst.out_buff_data[78] ;
 wire \top_inst.axis_out_inst.out_buff_data[79] ;
 wire \top_inst.axis_out_inst.out_buff_data[7] ;
 wire \top_inst.axis_out_inst.out_buff_data[80] ;
 wire \top_inst.axis_out_inst.out_buff_data[81] ;
 wire \top_inst.axis_out_inst.out_buff_data[82] ;
 wire \top_inst.axis_out_inst.out_buff_data[83] ;
 wire \top_inst.axis_out_inst.out_buff_data[84] ;
 wire \top_inst.axis_out_inst.out_buff_data[85] ;
 wire \top_inst.axis_out_inst.out_buff_data[86] ;
 wire \top_inst.axis_out_inst.out_buff_data[87] ;
 wire \top_inst.axis_out_inst.out_buff_data[88] ;
 wire \top_inst.axis_out_inst.out_buff_data[89] ;
 wire \top_inst.axis_out_inst.out_buff_data[8] ;
 wire \top_inst.axis_out_inst.out_buff_data[90] ;
 wire \top_inst.axis_out_inst.out_buff_data[91] ;
 wire \top_inst.axis_out_inst.out_buff_data[92] ;
 wire \top_inst.axis_out_inst.out_buff_data[93] ;
 wire \top_inst.axis_out_inst.out_buff_data[94] ;
 wire \top_inst.axis_out_inst.out_buff_data[95] ;
 wire \top_inst.axis_out_inst.out_buff_data[96] ;
 wire \top_inst.axis_out_inst.out_buff_data[97] ;
 wire \top_inst.axis_out_inst.out_buff_data[98] ;
 wire \top_inst.axis_out_inst.out_buff_data[99] ;
 wire \top_inst.axis_out_inst.out_buff_data[9] ;
 wire \top_inst.axis_out_inst.out_buff_enabled ;
 wire \top_inst.deskew_buff_inst.col_input[0] ;
 wire \top_inst.deskew_buff_inst.col_input[100] ;
 wire \top_inst.deskew_buff_inst.col_input[101] ;
 wire \top_inst.deskew_buff_inst.col_input[102] ;
 wire \top_inst.deskew_buff_inst.col_input[103] ;
 wire \top_inst.deskew_buff_inst.col_input[104] ;
 wire \top_inst.deskew_buff_inst.col_input[105] ;
 wire \top_inst.deskew_buff_inst.col_input[106] ;
 wire \top_inst.deskew_buff_inst.col_input[107] ;
 wire \top_inst.deskew_buff_inst.col_input[108] ;
 wire \top_inst.deskew_buff_inst.col_input[109] ;
 wire \top_inst.deskew_buff_inst.col_input[10] ;
 wire \top_inst.deskew_buff_inst.col_input[110] ;
 wire \top_inst.deskew_buff_inst.col_input[111] ;
 wire \top_inst.deskew_buff_inst.col_input[112] ;
 wire \top_inst.deskew_buff_inst.col_input[113] ;
 wire \top_inst.deskew_buff_inst.col_input[114] ;
 wire \top_inst.deskew_buff_inst.col_input[115] ;
 wire \top_inst.deskew_buff_inst.col_input[116] ;
 wire \top_inst.deskew_buff_inst.col_input[117] ;
 wire \top_inst.deskew_buff_inst.col_input[118] ;
 wire \top_inst.deskew_buff_inst.col_input[119] ;
 wire \top_inst.deskew_buff_inst.col_input[11] ;
 wire \top_inst.deskew_buff_inst.col_input[120] ;
 wire \top_inst.deskew_buff_inst.col_input[121] ;
 wire \top_inst.deskew_buff_inst.col_input[122] ;
 wire \top_inst.deskew_buff_inst.col_input[123] ;
 wire \top_inst.deskew_buff_inst.col_input[124] ;
 wire \top_inst.deskew_buff_inst.col_input[125] ;
 wire \top_inst.deskew_buff_inst.col_input[126] ;
 wire \top_inst.deskew_buff_inst.col_input[127] ;
 wire \top_inst.deskew_buff_inst.col_input[12] ;
 wire \top_inst.deskew_buff_inst.col_input[13] ;
 wire \top_inst.deskew_buff_inst.col_input[14] ;
 wire \top_inst.deskew_buff_inst.col_input[15] ;
 wire \top_inst.deskew_buff_inst.col_input[16] ;
 wire \top_inst.deskew_buff_inst.col_input[17] ;
 wire \top_inst.deskew_buff_inst.col_input[18] ;
 wire \top_inst.deskew_buff_inst.col_input[19] ;
 wire \top_inst.deskew_buff_inst.col_input[1] ;
 wire \top_inst.deskew_buff_inst.col_input[20] ;
 wire \top_inst.deskew_buff_inst.col_input[21] ;
 wire \top_inst.deskew_buff_inst.col_input[22] ;
 wire \top_inst.deskew_buff_inst.col_input[23] ;
 wire \top_inst.deskew_buff_inst.col_input[24] ;
 wire \top_inst.deskew_buff_inst.col_input[25] ;
 wire \top_inst.deskew_buff_inst.col_input[26] ;
 wire \top_inst.deskew_buff_inst.col_input[27] ;
 wire \top_inst.deskew_buff_inst.col_input[28] ;
 wire \top_inst.deskew_buff_inst.col_input[29] ;
 wire \top_inst.deskew_buff_inst.col_input[2] ;
 wire \top_inst.deskew_buff_inst.col_input[30] ;
 wire \top_inst.deskew_buff_inst.col_input[31] ;
 wire \top_inst.deskew_buff_inst.col_input[32] ;
 wire \top_inst.deskew_buff_inst.col_input[33] ;
 wire \top_inst.deskew_buff_inst.col_input[34] ;
 wire \top_inst.deskew_buff_inst.col_input[35] ;
 wire \top_inst.deskew_buff_inst.col_input[36] ;
 wire \top_inst.deskew_buff_inst.col_input[37] ;
 wire \top_inst.deskew_buff_inst.col_input[38] ;
 wire \top_inst.deskew_buff_inst.col_input[39] ;
 wire \top_inst.deskew_buff_inst.col_input[3] ;
 wire \top_inst.deskew_buff_inst.col_input[40] ;
 wire \top_inst.deskew_buff_inst.col_input[41] ;
 wire \top_inst.deskew_buff_inst.col_input[42] ;
 wire \top_inst.deskew_buff_inst.col_input[43] ;
 wire \top_inst.deskew_buff_inst.col_input[44] ;
 wire \top_inst.deskew_buff_inst.col_input[45] ;
 wire \top_inst.deskew_buff_inst.col_input[46] ;
 wire \top_inst.deskew_buff_inst.col_input[47] ;
 wire \top_inst.deskew_buff_inst.col_input[48] ;
 wire \top_inst.deskew_buff_inst.col_input[49] ;
 wire \top_inst.deskew_buff_inst.col_input[4] ;
 wire \top_inst.deskew_buff_inst.col_input[50] ;
 wire \top_inst.deskew_buff_inst.col_input[51] ;
 wire \top_inst.deskew_buff_inst.col_input[52] ;
 wire \top_inst.deskew_buff_inst.col_input[53] ;
 wire \top_inst.deskew_buff_inst.col_input[54] ;
 wire \top_inst.deskew_buff_inst.col_input[55] ;
 wire \top_inst.deskew_buff_inst.col_input[56] ;
 wire \top_inst.deskew_buff_inst.col_input[57] ;
 wire \top_inst.deskew_buff_inst.col_input[58] ;
 wire \top_inst.deskew_buff_inst.col_input[59] ;
 wire \top_inst.deskew_buff_inst.col_input[5] ;
 wire \top_inst.deskew_buff_inst.col_input[60] ;
 wire \top_inst.deskew_buff_inst.col_input[61] ;
 wire \top_inst.deskew_buff_inst.col_input[62] ;
 wire \top_inst.deskew_buff_inst.col_input[63] ;
 wire \top_inst.deskew_buff_inst.col_input[64] ;
 wire \top_inst.deskew_buff_inst.col_input[65] ;
 wire \top_inst.deskew_buff_inst.col_input[66] ;
 wire \top_inst.deskew_buff_inst.col_input[67] ;
 wire \top_inst.deskew_buff_inst.col_input[68] ;
 wire \top_inst.deskew_buff_inst.col_input[69] ;
 wire \top_inst.deskew_buff_inst.col_input[6] ;
 wire \top_inst.deskew_buff_inst.col_input[70] ;
 wire \top_inst.deskew_buff_inst.col_input[71] ;
 wire \top_inst.deskew_buff_inst.col_input[72] ;
 wire \top_inst.deskew_buff_inst.col_input[73] ;
 wire \top_inst.deskew_buff_inst.col_input[74] ;
 wire \top_inst.deskew_buff_inst.col_input[75] ;
 wire \top_inst.deskew_buff_inst.col_input[76] ;
 wire \top_inst.deskew_buff_inst.col_input[77] ;
 wire \top_inst.deskew_buff_inst.col_input[78] ;
 wire \top_inst.deskew_buff_inst.col_input[79] ;
 wire \top_inst.deskew_buff_inst.col_input[7] ;
 wire \top_inst.deskew_buff_inst.col_input[80] ;
 wire \top_inst.deskew_buff_inst.col_input[81] ;
 wire \top_inst.deskew_buff_inst.col_input[82] ;
 wire \top_inst.deskew_buff_inst.col_input[83] ;
 wire \top_inst.deskew_buff_inst.col_input[84] ;
 wire \top_inst.deskew_buff_inst.col_input[85] ;
 wire \top_inst.deskew_buff_inst.col_input[86] ;
 wire \top_inst.deskew_buff_inst.col_input[87] ;
 wire \top_inst.deskew_buff_inst.col_input[88] ;
 wire \top_inst.deskew_buff_inst.col_input[89] ;
 wire \top_inst.deskew_buff_inst.col_input[8] ;
 wire \top_inst.deskew_buff_inst.col_input[90] ;
 wire \top_inst.deskew_buff_inst.col_input[91] ;
 wire \top_inst.deskew_buff_inst.col_input[92] ;
 wire \top_inst.deskew_buff_inst.col_input[93] ;
 wire \top_inst.deskew_buff_inst.col_input[94] ;
 wire \top_inst.deskew_buff_inst.col_input[95] ;
 wire \top_inst.deskew_buff_inst.col_input[96] ;
 wire \top_inst.deskew_buff_inst.col_input[97] ;
 wire \top_inst.deskew_buff_inst.col_input[98] ;
 wire \top_inst.deskew_buff_inst.col_input[99] ;
 wire \top_inst.deskew_buff_inst.col_input[9] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][0] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][10] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][11] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][12] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][13] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][14] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][15] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][16] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][17] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][18] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][19] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][1] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][20] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][21] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][22] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][23] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][24] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][25] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][26] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][27] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][28] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][29] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][2] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][30] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][31] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][3] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][4] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][5] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][6] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][7] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][8] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][9] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][0] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][10] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][11] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][12] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][13] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][14] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][15] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][16] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][17] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][18] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][19] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][1] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][20] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][21] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][22] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][23] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][24] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][25] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][26] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][27] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][28] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][29] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][2] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][30] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][31] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][3] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][4] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][5] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][6] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][7] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][8] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][9] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][0] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][10] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][11] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][12] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][13] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][14] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][15] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][16] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][17] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][18] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][19] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][1] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][20] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][21] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][22] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][23] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][24] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][25] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][26] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][27] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][28] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][29] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][2] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][30] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][31] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][3] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][4] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][5] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][6] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][7] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][8] ;
 wire \top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][9] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][0] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][10] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][11] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][12] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][13] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][14] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][15] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][16] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][17] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][18] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][19] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][1] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][20] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][21] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][22] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][23] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][24] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][25] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][26] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][27] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][28] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][29] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][2] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][30] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][31] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][3] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][4] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][5] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][6] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][7] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][8] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][9] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][0] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][10] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][11] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][12] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][13] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][14] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][15] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][16] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][17] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][18] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][19] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][1] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][20] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][21] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][22] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][23] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][24] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][25] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][26] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][27] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][28] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][29] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][2] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][30] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][31] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][3] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][4] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][5] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][6] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][7] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][8] ;
 wire \top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][9] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][0] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][10] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][11] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][12] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][13] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][14] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][15] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][16] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][17] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][18] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][19] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][1] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][20] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][21] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][22] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][23] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][24] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][25] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][26] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][27] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][28] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][29] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][2] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][30] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][31] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][3] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][4] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][5] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][6] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][7] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][8] ;
 wire \top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][9] ;
 wire \top_inst.grid_inst.data_path_wires[11][0] ;
 wire \top_inst.grid_inst.data_path_wires[11][1] ;
 wire \top_inst.grid_inst.data_path_wires[11][2] ;
 wire \top_inst.grid_inst.data_path_wires[11][3] ;
 wire \top_inst.grid_inst.data_path_wires[11][4] ;
 wire \top_inst.grid_inst.data_path_wires[11][5] ;
 wire \top_inst.grid_inst.data_path_wires[11][6] ;
 wire \top_inst.grid_inst.data_path_wires[11][7] ;
 wire \top_inst.grid_inst.data_path_wires[12][0] ;
 wire \top_inst.grid_inst.data_path_wires[12][1] ;
 wire \top_inst.grid_inst.data_path_wires[12][2] ;
 wire \top_inst.grid_inst.data_path_wires[12][3] ;
 wire \top_inst.grid_inst.data_path_wires[12][4] ;
 wire \top_inst.grid_inst.data_path_wires[12][5] ;
 wire \top_inst.grid_inst.data_path_wires[12][6] ;
 wire \top_inst.grid_inst.data_path_wires[12][7] ;
 wire \top_inst.grid_inst.data_path_wires[13][0] ;
 wire \top_inst.grid_inst.data_path_wires[13][1] ;
 wire \top_inst.grid_inst.data_path_wires[13][2] ;
 wire \top_inst.grid_inst.data_path_wires[13][3] ;
 wire \top_inst.grid_inst.data_path_wires[13][4] ;
 wire \top_inst.grid_inst.data_path_wires[13][5] ;
 wire \top_inst.grid_inst.data_path_wires[13][6] ;
 wire \top_inst.grid_inst.data_path_wires[13][7] ;
 wire \top_inst.grid_inst.data_path_wires[16][0] ;
 wire \top_inst.grid_inst.data_path_wires[16][1] ;
 wire \top_inst.grid_inst.data_path_wires[16][2] ;
 wire \top_inst.grid_inst.data_path_wires[16][3] ;
 wire \top_inst.grid_inst.data_path_wires[16][4] ;
 wire \top_inst.grid_inst.data_path_wires[16][5] ;
 wire \top_inst.grid_inst.data_path_wires[16][6] ;
 wire \top_inst.grid_inst.data_path_wires[16][7] ;
 wire \top_inst.grid_inst.data_path_wires[17][0] ;
 wire \top_inst.grid_inst.data_path_wires[17][1] ;
 wire \top_inst.grid_inst.data_path_wires[17][2] ;
 wire \top_inst.grid_inst.data_path_wires[17][3] ;
 wire \top_inst.grid_inst.data_path_wires[17][4] ;
 wire \top_inst.grid_inst.data_path_wires[17][5] ;
 wire \top_inst.grid_inst.data_path_wires[17][6] ;
 wire \top_inst.grid_inst.data_path_wires[17][7] ;
 wire \top_inst.grid_inst.data_path_wires[18][0] ;
 wire \top_inst.grid_inst.data_path_wires[18][1] ;
 wire \top_inst.grid_inst.data_path_wires[18][2] ;
 wire \top_inst.grid_inst.data_path_wires[18][3] ;
 wire \top_inst.grid_inst.data_path_wires[18][4] ;
 wire \top_inst.grid_inst.data_path_wires[18][5] ;
 wire \top_inst.grid_inst.data_path_wires[18][6] ;
 wire \top_inst.grid_inst.data_path_wires[18][7] ;
 wire \top_inst.grid_inst.data_path_wires[1][0] ;
 wire \top_inst.grid_inst.data_path_wires[1][1] ;
 wire \top_inst.grid_inst.data_path_wires[1][2] ;
 wire \top_inst.grid_inst.data_path_wires[1][3] ;
 wire \top_inst.grid_inst.data_path_wires[1][4] ;
 wire \top_inst.grid_inst.data_path_wires[1][5] ;
 wire \top_inst.grid_inst.data_path_wires[1][6] ;
 wire \top_inst.grid_inst.data_path_wires[1][7] ;
 wire \top_inst.grid_inst.data_path_wires[2][0] ;
 wire \top_inst.grid_inst.data_path_wires[2][1] ;
 wire \top_inst.grid_inst.data_path_wires[2][2] ;
 wire \top_inst.grid_inst.data_path_wires[2][3] ;
 wire \top_inst.grid_inst.data_path_wires[2][4] ;
 wire \top_inst.grid_inst.data_path_wires[2][5] ;
 wire \top_inst.grid_inst.data_path_wires[2][6] ;
 wire \top_inst.grid_inst.data_path_wires[2][7] ;
 wire \top_inst.grid_inst.data_path_wires[3][0] ;
 wire \top_inst.grid_inst.data_path_wires[3][1] ;
 wire \top_inst.grid_inst.data_path_wires[3][2] ;
 wire \top_inst.grid_inst.data_path_wires[3][3] ;
 wire \top_inst.grid_inst.data_path_wires[3][4] ;
 wire \top_inst.grid_inst.data_path_wires[3][5] ;
 wire \top_inst.grid_inst.data_path_wires[3][6] ;
 wire \top_inst.grid_inst.data_path_wires[3][7] ;
 wire \top_inst.grid_inst.data_path_wires[6][0] ;
 wire \top_inst.grid_inst.data_path_wires[6][1] ;
 wire \top_inst.grid_inst.data_path_wires[6][2] ;
 wire \top_inst.grid_inst.data_path_wires[6][3] ;
 wire \top_inst.grid_inst.data_path_wires[6][4] ;
 wire \top_inst.grid_inst.data_path_wires[6][5] ;
 wire \top_inst.grid_inst.data_path_wires[6][6] ;
 wire \top_inst.grid_inst.data_path_wires[6][7] ;
 wire \top_inst.grid_inst.data_path_wires[7][0] ;
 wire \top_inst.grid_inst.data_path_wires[7][1] ;
 wire \top_inst.grid_inst.data_path_wires[7][2] ;
 wire \top_inst.grid_inst.data_path_wires[7][3] ;
 wire \top_inst.grid_inst.data_path_wires[7][4] ;
 wire \top_inst.grid_inst.data_path_wires[7][5] ;
 wire \top_inst.grid_inst.data_path_wires[7][6] ;
 wire \top_inst.grid_inst.data_path_wires[7][7] ;
 wire \top_inst.grid_inst.data_path_wires[8][0] ;
 wire \top_inst.grid_inst.data_path_wires[8][1] ;
 wire \top_inst.grid_inst.data_path_wires[8][2] ;
 wire \top_inst.grid_inst.data_path_wires[8][3] ;
 wire \top_inst.grid_inst.data_path_wires[8][4] ;
 wire \top_inst.grid_inst.data_path_wires[8][5] ;
 wire \top_inst.grid_inst.data_path_wires[8][6] ;
 wire \top_inst.grid_inst.data_path_wires[8][7] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[0] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[10] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[11] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[12] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[13] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[14] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[15] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[1] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[2] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[3] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[4] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[5] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[6] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[7] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[8] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[9] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[7] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[0] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[10] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[11] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[12] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[13] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[14] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[15] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[1] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[2] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[3] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[4] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[5] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[6] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[7] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[8] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[9] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[7] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[0] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[10] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[11] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[12] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[13] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[14] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[15] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[1] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[2] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[3] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[4] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[5] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[6] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[7] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[8] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[9] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[7] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[0] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[10] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[11] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[12] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[13] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[14] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[15] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[1] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[2] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[3] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[4] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[5] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[6] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[7] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[8] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[9] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[7] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[0] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[10] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[11] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[12] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[13] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[14] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[15] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[16] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[17] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[18] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[19] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[1] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[20] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[21] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[23] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[24] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[25] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[27] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[2] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[31] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[3] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[4] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[5] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[6] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[7] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[8] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[9] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[7] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[0] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[10] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[11] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[12] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[13] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[14] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[15] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[16] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[1] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[2] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[3] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[4] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[5] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[6] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[7] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[8] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[9] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[7] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[0] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[10] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[11] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[12] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[13] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[14] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[15] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[16] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[1] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[2] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[3] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[4] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[5] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[6] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[7] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[8] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[9] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[7] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[0] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[10] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[11] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[12] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[13] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[14] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[15] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[16] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[1] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[2] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[3] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[4] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[5] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[6] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[7] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[8] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[9] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[7] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[0] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[10] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[11] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[12] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[13] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[14] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[15] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[16] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[17] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[18] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[19] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[1] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[20] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[21] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[22] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[23] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[24] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[25] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[26] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[27] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[28] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[29] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[2] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[30] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[31] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[3] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[4] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[5] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[6] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[7] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[8] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[9] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[7] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[0] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[10] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[11] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[12] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[13] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[14] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[15] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[16] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[17] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[18] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[19] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[1] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[20] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[21] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[23] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[24] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[25] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[27] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[2] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[31] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[3] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[4] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[5] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[6] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[7] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[8] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[9] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[7] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[0] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[10] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[11] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[12] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[13] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[14] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[15] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[16] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[17] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[18] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[19] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[1] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[20] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[21] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[23] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[24] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[25] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[27] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[2] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[31] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[3] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[4] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[5] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[6] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[7] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[8] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[9] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[7] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[0] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[10] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[11] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[12] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[13] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[14] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[15] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[16] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[17] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[18] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[19] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[1] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[20] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[21] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[23] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[24] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[25] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[27] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[2] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[31] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[3] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[4] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[5] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[6] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[7] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[8] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[9] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[7] ;
 wire \top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[7] ;
 wire \top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[7] ;
 wire \top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[7] ;
 wire \top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[0] ;
 wire \top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[1] ;
 wire \top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[2] ;
 wire \top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[3] ;
 wire \top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[4] ;
 wire \top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[5] ;
 wire \top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[6] ;
 wire \top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[7] ;
 wire \top_inst.skew_buff_inst.row[0].output_reg[0] ;
 wire \top_inst.skew_buff_inst.row[0].output_reg[1] ;
 wire \top_inst.skew_buff_inst.row[0].output_reg[2] ;
 wire \top_inst.skew_buff_inst.row[0].output_reg[3] ;
 wire \top_inst.skew_buff_inst.row[0].output_reg[4] ;
 wire \top_inst.skew_buff_inst.row[0].output_reg[5] ;
 wire \top_inst.skew_buff_inst.row[0].output_reg[6] ;
 wire \top_inst.skew_buff_inst.row[0].output_reg[7] ;
 wire \top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][0] ;
 wire \top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][1] ;
 wire \top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][2] ;
 wire \top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][3] ;
 wire \top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][4] ;
 wire \top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][5] ;
 wire \top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][6] ;
 wire \top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][7] ;
 wire \top_inst.skew_buff_inst.row[1].output_reg[0] ;
 wire \top_inst.skew_buff_inst.row[1].output_reg[1] ;
 wire \top_inst.skew_buff_inst.row[1].output_reg[2] ;
 wire \top_inst.skew_buff_inst.row[1].output_reg[3] ;
 wire \top_inst.skew_buff_inst.row[1].output_reg[4] ;
 wire \top_inst.skew_buff_inst.row[1].output_reg[5] ;
 wire \top_inst.skew_buff_inst.row[1].output_reg[6] ;
 wire \top_inst.skew_buff_inst.row[1].output_reg[7] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][0] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][1] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][2] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][3] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][4] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][5] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][6] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][7] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][0] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][1] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][2] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][3] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][4] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][5] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][6] ;
 wire \top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][7] ;
 wire \top_inst.skew_buff_inst.row[2].output_reg[0] ;
 wire \top_inst.skew_buff_inst.row[2].output_reg[1] ;
 wire \top_inst.skew_buff_inst.row[2].output_reg[2] ;
 wire \top_inst.skew_buff_inst.row[2].output_reg[3] ;
 wire \top_inst.skew_buff_inst.row[2].output_reg[4] ;
 wire \top_inst.skew_buff_inst.row[2].output_reg[5] ;
 wire \top_inst.skew_buff_inst.row[2].output_reg[6] ;
 wire \top_inst.skew_buff_inst.row[2].output_reg[7] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][0] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][1] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][2] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][3] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][4] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][5] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][6] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][7] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][0] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][1] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][2] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][3] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][4] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][5] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][6] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][7] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][0] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][1] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][2] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][3] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][4] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][5] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][6] ;
 wire \top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][7] ;
 wire \top_inst.skew_buff_inst.row[3].output_reg[0] ;
 wire \top_inst.skew_buff_inst.row[3].output_reg[1] ;
 wire \top_inst.skew_buff_inst.row[3].output_reg[2] ;
 wire \top_inst.skew_buff_inst.row[3].output_reg[3] ;
 wire \top_inst.skew_buff_inst.row[3].output_reg[4] ;
 wire \top_inst.skew_buff_inst.row[3].output_reg[5] ;
 wire \top_inst.skew_buff_inst.row[3].output_reg[6] ;
 wire \top_inst.skew_buff_inst.row[3].output_reg[7] ;
 wire \top_inst.valid_pipe[0] ;
 wire \top_inst.valid_pipe[1] ;
 wire \top_inst.valid_pipe[2] ;
 wire \top_inst.valid_pipe[3] ;
 wire \top_inst.valid_pipe[4] ;
 wire \top_inst.valid_pipe[5] ;
 wire \top_inst.valid_pipe[6] ;
 wire \top_inst.valid_pipe[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_4_0__leaf_clk;
 wire clknet_4_1__leaf_clk;
 wire clknet_4_2__leaf_clk;
 wire clknet_4_3__leaf_clk;
 wire clknet_4_4__leaf_clk;
 wire clknet_4_5__leaf_clk;
 wire clknet_4_6__leaf_clk;
 wire clknet_4_7__leaf_clk;
 wire clknet_4_8__leaf_clk;
 wire clknet_4_9__leaf_clk;
 wire clknet_4_10__leaf_clk;
 wire clknet_4_11__leaf_clk;
 wire clknet_4_12__leaf_clk;
 wire clknet_4_13__leaf_clk;
 wire clknet_4_14__leaf_clk;
 wire clknet_4_15__leaf_clk;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net252;
 wire net253;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;

 sky130_fd_sc_hd__nor2b_4 _11733_ (.A(net35),
    .B_N(net166),
    .Y(_04856_));
 sky130_fd_sc_hd__nand2_8 _11734_ (.A(\top_inst.axis_in_inst.inbuf_valid ),
    .B(_04856_),
    .Y(net37));
 sky130_fd_sc_hd__nand2b_4 _11735_ (.A_N(net35),
    .B(net166),
    .Y(_04857_));
 sky130_fd_sc_hd__nand2_8 _11736_ (.A(\top_inst.axis_in_inst.inbuf_valid ),
    .B(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__buf_8 _11737_ (.A(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__buf_4 _11738_ (.A(_04859_),
    .X(_04860_));
 sky130_fd_sc_hd__inv_6 _11739_ (.A(\top_inst.axis_in_inst.inbuf_valid ),
    .Y(_04861_));
 sky130_fd_sc_hd__nor2_1 _11740_ (.A(_04861_),
    .B(_04856_),
    .Y(_04862_));
 sky130_fd_sc_hd__buf_8 _11741_ (.A(_04862_),
    .X(_04863_));
 sky130_fd_sc_hd__buf_2 _11742_ (.A(_04863_),
    .X(_04864_));
 sky130_fd_sc_hd__buf_4 _11743_ (.A(_04864_),
    .X(_04865_));
 sky130_fd_sc_hd__or2_1 _11744_ (.A(\top_inst.axis_out_inst.out_buff_data[121] ),
    .B(_04865_),
    .X(_04866_));
 sky130_fd_sc_hd__buf_8 _11745_ (.A(net36),
    .X(_04867_));
 sky130_fd_sc_hd__inv_2 _11746_ (.A(_04867_),
    .Y(_04868_));
 sky130_fd_sc_hd__clkbuf_8 _11747_ (.A(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__buf_8 _11748_ (.A(_04869_),
    .X(_04870_));
 sky130_fd_sc_hd__o211a_1 _11749_ (.A1(net777),
    .A2(_04860_),
    .B1(_04866_),
    .C1(_04870_),
    .X(_00000_));
 sky130_fd_sc_hd__or2_1 _11750_ (.A(net451),
    .B(_04865_),
    .X(_04871_));
 sky130_fd_sc_hd__o211a_1 _11751_ (.A1(net630),
    .A2(_04860_),
    .B1(_04871_),
    .C1(_04870_),
    .X(_00001_));
 sky130_fd_sc_hd__or2_1 _11752_ (.A(net410),
    .B(_04865_),
    .X(_04872_));
 sky130_fd_sc_hd__buf_6 _11753_ (.A(_04868_),
    .X(_04873_));
 sky130_fd_sc_hd__buf_4 _11754_ (.A(_04873_),
    .X(_04874_));
 sky130_fd_sc_hd__buf_4 _11755_ (.A(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__o211a_1 _11756_ (.A1(net724),
    .A2(_04860_),
    .B1(_04872_),
    .C1(_04875_),
    .X(_00002_));
 sky130_fd_sc_hd__clkbuf_4 _11757_ (.A(_04863_),
    .X(_04876_));
 sky130_fd_sc_hd__buf_4 _11758_ (.A(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__or2_1 _11759_ (.A(\top_inst.axis_out_inst.out_buff_data[124] ),
    .B(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__o211a_1 _11760_ (.A1(net564),
    .A2(_04860_),
    .B1(_04878_),
    .C1(_04875_),
    .X(_00003_));
 sky130_fd_sc_hd__or2_1 _11761_ (.A(\top_inst.axis_out_inst.out_buff_data[125] ),
    .B(_04877_),
    .X(_04879_));
 sky130_fd_sc_hd__o211a_1 _11762_ (.A1(net666),
    .A2(_04860_),
    .B1(_04879_),
    .C1(_04875_),
    .X(_00004_));
 sky130_fd_sc_hd__or2_1 _11763_ (.A(\top_inst.axis_out_inst.out_buff_data[126] ),
    .B(_04877_),
    .X(_04880_));
 sky130_fd_sc_hd__o211a_1 _11764_ (.A1(net471),
    .A2(_04860_),
    .B1(_04880_),
    .C1(_04875_),
    .X(_00005_));
 sky130_fd_sc_hd__or2_1 _11765_ (.A(\top_inst.axis_out_inst.out_buff_data[127] ),
    .B(_04877_),
    .X(_04881_));
 sky130_fd_sc_hd__o211a_1 _11766_ (.A1(net499),
    .A2(_04860_),
    .B1(_04881_),
    .C1(_04875_),
    .X(_00006_));
 sky130_fd_sc_hd__or2_1 _11767_ (.A(\top_inst.axis_out_inst.out_buff_data[64] ),
    .B(_04877_),
    .X(_04882_));
 sky130_fd_sc_hd__o211a_1 _11768_ (.A1(net625),
    .A2(_04860_),
    .B1(_04882_),
    .C1(_04875_),
    .X(_00007_));
 sky130_fd_sc_hd__or2_1 _11769_ (.A(net622),
    .B(_04877_),
    .X(_04883_));
 sky130_fd_sc_hd__o211a_1 _11770_ (.A1(net744),
    .A2(_04860_),
    .B1(_04883_),
    .C1(_04875_),
    .X(_00008_));
 sky130_fd_sc_hd__or2_1 _11771_ (.A(net364),
    .B(_04877_),
    .X(_04884_));
 sky130_fd_sc_hd__o211a_1 _11772_ (.A1(net888),
    .A2(_04860_),
    .B1(_04884_),
    .C1(_04875_),
    .X(_00009_));
 sky130_fd_sc_hd__clkbuf_4 _11773_ (.A(_04859_),
    .X(_04885_));
 sky130_fd_sc_hd__or2_1 _11774_ (.A(net377),
    .B(_04877_),
    .X(_04886_));
 sky130_fd_sc_hd__o211a_1 _11775_ (.A1(net594),
    .A2(_04885_),
    .B1(_04886_),
    .C1(_04875_),
    .X(_00010_));
 sky130_fd_sc_hd__or2_1 _11776_ (.A(\top_inst.axis_out_inst.out_buff_data[68] ),
    .B(_04877_),
    .X(_04887_));
 sky130_fd_sc_hd__o211a_1 _11777_ (.A1(net348),
    .A2(_04885_),
    .B1(_04887_),
    .C1(_04875_),
    .X(_00011_));
 sky130_fd_sc_hd__or2_1 _11778_ (.A(\top_inst.axis_out_inst.out_buff_data[69] ),
    .B(_04877_),
    .X(_04888_));
 sky130_fd_sc_hd__buf_2 _11779_ (.A(_04874_),
    .X(_04889_));
 sky130_fd_sc_hd__o211a_1 _11780_ (.A1(net362),
    .A2(_04885_),
    .B1(_04888_),
    .C1(_04889_),
    .X(_00012_));
 sky130_fd_sc_hd__buf_2 _11781_ (.A(_04876_),
    .X(_04890_));
 sky130_fd_sc_hd__or2_1 _11782_ (.A(\top_inst.axis_out_inst.out_buff_data[70] ),
    .B(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__o211a_1 _11783_ (.A1(net360),
    .A2(_04885_),
    .B1(_04891_),
    .C1(_04889_),
    .X(_00013_));
 sky130_fd_sc_hd__or2_1 _11784_ (.A(\top_inst.axis_out_inst.out_buff_data[71] ),
    .B(_04890_),
    .X(_04892_));
 sky130_fd_sc_hd__o211a_1 _11785_ (.A1(net337),
    .A2(_04885_),
    .B1(_04892_),
    .C1(_04889_),
    .X(_00014_));
 sky130_fd_sc_hd__or2_1 _11786_ (.A(net757),
    .B(_04890_),
    .X(_04893_));
 sky130_fd_sc_hd__o211a_1 _11787_ (.A1(net803),
    .A2(_04885_),
    .B1(_04893_),
    .C1(_04889_),
    .X(_00015_));
 sky130_fd_sc_hd__or2_1 _11788_ (.A(\top_inst.axis_out_inst.out_buff_data[73] ),
    .B(_04890_),
    .X(_04894_));
 sky130_fd_sc_hd__o211a_1 _11789_ (.A1(net367),
    .A2(_04885_),
    .B1(_04894_),
    .C1(_04889_),
    .X(_00016_));
 sky130_fd_sc_hd__or2_1 _11790_ (.A(net743),
    .B(_04890_),
    .X(_04895_));
 sky130_fd_sc_hd__o211a_1 _11791_ (.A1(net866),
    .A2(_04885_),
    .B1(_04895_),
    .C1(_04889_),
    .X(_00017_));
 sky130_fd_sc_hd__or2_1 _11792_ (.A(net727),
    .B(_04890_),
    .X(_04896_));
 sky130_fd_sc_hd__o211a_1 _11793_ (.A1(net829),
    .A2(_04885_),
    .B1(_04896_),
    .C1(_04889_),
    .X(_00018_));
 sky130_fd_sc_hd__or2_1 _11794_ (.A(net705),
    .B(_04890_),
    .X(_04897_));
 sky130_fd_sc_hd__o211a_1 _11795_ (.A1(net857),
    .A2(_04885_),
    .B1(_04897_),
    .C1(_04889_),
    .X(_00019_));
 sky130_fd_sc_hd__clkbuf_4 _11796_ (.A(_04859_),
    .X(_04898_));
 sky130_fd_sc_hd__or2_1 _11797_ (.A(net468),
    .B(_04890_),
    .X(_04899_));
 sky130_fd_sc_hd__o211a_1 _11798_ (.A1(net856),
    .A2(_04898_),
    .B1(_04899_),
    .C1(_04889_),
    .X(_00020_));
 sky130_fd_sc_hd__or2_1 _11799_ (.A(\top_inst.axis_out_inst.out_buff_data[78] ),
    .B(_04890_),
    .X(_04900_));
 sky130_fd_sc_hd__o211a_1 _11800_ (.A1(net570),
    .A2(_04898_),
    .B1(_04900_),
    .C1(_04889_),
    .X(_00021_));
 sky130_fd_sc_hd__or2_1 _11801_ (.A(\top_inst.axis_out_inst.out_buff_data[79] ),
    .B(_04890_),
    .X(_04901_));
 sky130_fd_sc_hd__clkbuf_4 _11802_ (.A(_04874_),
    .X(_04902_));
 sky130_fd_sc_hd__o211a_1 _11803_ (.A1(net614),
    .A2(_04898_),
    .B1(_04901_),
    .C1(_04902_),
    .X(_00022_));
 sky130_fd_sc_hd__buf_2 _11804_ (.A(_04876_),
    .X(_04903_));
 sky130_fd_sc_hd__or2_1 _11805_ (.A(\top_inst.axis_out_inst.out_buff_data[80] ),
    .B(_04903_),
    .X(_04904_));
 sky130_fd_sc_hd__o211a_1 _11806_ (.A1(net640),
    .A2(_04898_),
    .B1(_04904_),
    .C1(_04902_),
    .X(_00023_));
 sky130_fd_sc_hd__or2_1 _11807_ (.A(net462),
    .B(_04903_),
    .X(_04905_));
 sky130_fd_sc_hd__o211a_1 _11808_ (.A1(net576),
    .A2(_04898_),
    .B1(_04905_),
    .C1(_04902_),
    .X(_00024_));
 sky130_fd_sc_hd__or2_1 _11809_ (.A(\top_inst.axis_out_inst.out_buff_data[82] ),
    .B(_04903_),
    .X(_04906_));
 sky130_fd_sc_hd__o211a_1 _11810_ (.A1(net522),
    .A2(_04898_),
    .B1(_04906_),
    .C1(_04902_),
    .X(_00025_));
 sky130_fd_sc_hd__or2_1 _11811_ (.A(net742),
    .B(_04903_),
    .X(_04907_));
 sky130_fd_sc_hd__o211a_1 _11812_ (.A1(net800),
    .A2(_04898_),
    .B1(_04907_),
    .C1(_04902_),
    .X(_00026_));
 sky130_fd_sc_hd__or2_1 _11813_ (.A(net393),
    .B(_04903_),
    .X(_04908_));
 sky130_fd_sc_hd__o211a_1 _11814_ (.A1(net933),
    .A2(_04898_),
    .B1(_04908_),
    .C1(_04902_),
    .X(_00027_));
 sky130_fd_sc_hd__or2_1 _11815_ (.A(net391),
    .B(_04903_),
    .X(_04909_));
 sky130_fd_sc_hd__o211a_1 _11816_ (.A1(net908),
    .A2(_04898_),
    .B1(_04909_),
    .C1(_04902_),
    .X(_00028_));
 sky130_fd_sc_hd__or2_1 _11817_ (.A(\top_inst.axis_out_inst.out_buff_data[86] ),
    .B(_04903_),
    .X(_04910_));
 sky130_fd_sc_hd__o211a_1 _11818_ (.A1(net474),
    .A2(_04898_),
    .B1(_04910_),
    .C1(_04902_),
    .X(_00029_));
 sky130_fd_sc_hd__buf_4 _11819_ (.A(_04858_),
    .X(_04911_));
 sky130_fd_sc_hd__clkbuf_4 _11820_ (.A(_04911_),
    .X(_04912_));
 sky130_fd_sc_hd__or2_1 _11821_ (.A(net629),
    .B(_04903_),
    .X(_04913_));
 sky130_fd_sc_hd__o211a_1 _11822_ (.A1(net865),
    .A2(_04912_),
    .B1(_04913_),
    .C1(_04902_),
    .X(_00030_));
 sky130_fd_sc_hd__or2_1 _11823_ (.A(net657),
    .B(_04903_),
    .X(_04914_));
 sky130_fd_sc_hd__o211a_1 _11824_ (.A1(net889),
    .A2(_04912_),
    .B1(_04914_),
    .C1(_04902_),
    .X(_00031_));
 sky130_fd_sc_hd__or2_1 _11825_ (.A(net415),
    .B(_04903_),
    .X(_04915_));
 sky130_fd_sc_hd__clkbuf_4 _11826_ (.A(_04874_),
    .X(_04916_));
 sky130_fd_sc_hd__o211a_1 _11827_ (.A1(net652),
    .A2(_04912_),
    .B1(_04915_),
    .C1(_04916_),
    .X(_00032_));
 sky130_fd_sc_hd__buf_2 _11828_ (.A(_04876_),
    .X(_04917_));
 sky130_fd_sc_hd__or2_1 _11829_ (.A(net694),
    .B(_04917_),
    .X(_04918_));
 sky130_fd_sc_hd__o211a_1 _11830_ (.A1(net794),
    .A2(_04912_),
    .B1(_04918_),
    .C1(_04916_),
    .X(_00033_));
 sky130_fd_sc_hd__or2_1 _11831_ (.A(net599),
    .B(_04917_),
    .X(_04919_));
 sky130_fd_sc_hd__o211a_1 _11832_ (.A1(net688),
    .A2(_04912_),
    .B1(_04919_),
    .C1(_04916_),
    .X(_00034_));
 sky130_fd_sc_hd__or2_1 _11833_ (.A(net434),
    .B(_04917_),
    .X(_04920_));
 sky130_fd_sc_hd__o211a_1 _11834_ (.A1(net944),
    .A2(_04912_),
    .B1(_04920_),
    .C1(_04916_),
    .X(_00035_));
 sky130_fd_sc_hd__or2_1 _11835_ (.A(\top_inst.axis_out_inst.out_buff_data[93] ),
    .B(_04917_),
    .X(_04921_));
 sky130_fd_sc_hd__o211a_1 _11836_ (.A1(net684),
    .A2(_04912_),
    .B1(_04921_),
    .C1(_04916_),
    .X(_00036_));
 sky130_fd_sc_hd__or2_1 _11837_ (.A(\top_inst.axis_out_inst.out_buff_data[94] ),
    .B(_04917_),
    .X(_04922_));
 sky130_fd_sc_hd__o211a_1 _11838_ (.A1(net689),
    .A2(_04912_),
    .B1(_04922_),
    .C1(_04916_),
    .X(_00037_));
 sky130_fd_sc_hd__or2_1 _11839_ (.A(\top_inst.axis_out_inst.out_buff_data[95] ),
    .B(_04917_),
    .X(_04923_));
 sky130_fd_sc_hd__o211a_1 _11840_ (.A1(net428),
    .A2(_04912_),
    .B1(_04923_),
    .C1(_04916_),
    .X(_00038_));
 sky130_fd_sc_hd__or2_1 _11841_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][0] ),
    .B(_04917_),
    .X(_04924_));
 sky130_fd_sc_hd__o211a_1 _11842_ (.A1(net454),
    .A2(_04912_),
    .B1(_04924_),
    .C1(_04916_),
    .X(_00039_));
 sky130_fd_sc_hd__clkbuf_4 _11843_ (.A(_04911_),
    .X(_04925_));
 sky130_fd_sc_hd__or2_1 _11844_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][1] ),
    .B(_04917_),
    .X(_04926_));
 sky130_fd_sc_hd__o211a_1 _11845_ (.A1(net325),
    .A2(_04925_),
    .B1(_04926_),
    .C1(_04916_),
    .X(_00040_));
 sky130_fd_sc_hd__or2_1 _11846_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][2] ),
    .B(_04917_),
    .X(_04927_));
 sky130_fd_sc_hd__o211a_1 _11847_ (.A1(net282),
    .A2(_04925_),
    .B1(_04927_),
    .C1(_04916_),
    .X(_00041_));
 sky130_fd_sc_hd__or2_1 _11848_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][3] ),
    .B(_04917_),
    .X(_04928_));
 sky130_fd_sc_hd__buf_2 _11849_ (.A(_04874_),
    .X(_04929_));
 sky130_fd_sc_hd__o211a_1 _11850_ (.A1(net313),
    .A2(_04925_),
    .B1(_04928_),
    .C1(_04929_),
    .X(_00042_));
 sky130_fd_sc_hd__clkbuf_2 _11851_ (.A(_04876_),
    .X(_04930_));
 sky130_fd_sc_hd__or2_1 _11852_ (.A(net348),
    .B(_04930_),
    .X(_04931_));
 sky130_fd_sc_hd__o211a_1 _11853_ (.A1(net604),
    .A2(_04925_),
    .B1(_04931_),
    .C1(_04929_),
    .X(_00043_));
 sky130_fd_sc_hd__or2_1 _11854_ (.A(net362),
    .B(_04930_),
    .X(_04932_));
 sky130_fd_sc_hd__o211a_1 _11855_ (.A1(net921),
    .A2(_04925_),
    .B1(_04932_),
    .C1(_04929_),
    .X(_00044_));
 sky130_fd_sc_hd__or2_1 _11856_ (.A(net360),
    .B(_04930_),
    .X(_04933_));
 sky130_fd_sc_hd__o211a_1 _11857_ (.A1(net860),
    .A2(_04925_),
    .B1(_04933_),
    .C1(_04929_),
    .X(_00045_));
 sky130_fd_sc_hd__or2_1 _11858_ (.A(net337),
    .B(_04930_),
    .X(_04934_));
 sky130_fd_sc_hd__o211a_1 _11859_ (.A1(net938),
    .A2(_04925_),
    .B1(_04934_),
    .C1(_04929_),
    .X(_00046_));
 sky130_fd_sc_hd__or2_1 _11860_ (.A(net803),
    .B(_04930_),
    .X(_04935_));
 sky130_fd_sc_hd__o211a_1 _11861_ (.A1(net808),
    .A2(_04925_),
    .B1(_04935_),
    .C1(_04929_),
    .X(_00047_));
 sky130_fd_sc_hd__or2_1 _11862_ (.A(net367),
    .B(_04930_),
    .X(_04936_));
 sky130_fd_sc_hd__o211a_1 _11863_ (.A1(net924),
    .A2(_04925_),
    .B1(_04936_),
    .C1(_04929_),
    .X(_00048_));
 sky130_fd_sc_hd__or2_1 _11864_ (.A(net866),
    .B(_04930_),
    .X(_04937_));
 sky130_fd_sc_hd__o211a_1 _11865_ (.A1(net897),
    .A2(_04925_),
    .B1(_04937_),
    .C1(_04929_),
    .X(_00049_));
 sky130_fd_sc_hd__clkbuf_4 _11866_ (.A(_04911_),
    .X(_04938_));
 sky130_fd_sc_hd__or2_1 _11867_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][11] ),
    .B(_04930_),
    .X(_04939_));
 sky130_fd_sc_hd__o211a_1 _11868_ (.A1(net753),
    .A2(_04938_),
    .B1(_04939_),
    .C1(_04929_),
    .X(_00050_));
 sky130_fd_sc_hd__or2_1 _11869_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][12] ),
    .B(_04930_),
    .X(_04940_));
 sky130_fd_sc_hd__o211a_1 _11870_ (.A1(net839),
    .A2(_04938_),
    .B1(_04940_),
    .C1(_04929_),
    .X(_00051_));
 sky130_fd_sc_hd__or2_1 _11871_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][13] ),
    .B(_04930_),
    .X(_04941_));
 sky130_fd_sc_hd__buf_2 _11872_ (.A(_04874_),
    .X(_04942_));
 sky130_fd_sc_hd__o211a_1 _11873_ (.A1(net818),
    .A2(_04938_),
    .B1(_04941_),
    .C1(_04942_),
    .X(_00052_));
 sky130_fd_sc_hd__buf_2 _11874_ (.A(_04876_),
    .X(_04943_));
 sky130_fd_sc_hd__or2_1 _11875_ (.A(net570),
    .B(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__o211a_1 _11876_ (.A1(net611),
    .A2(_04938_),
    .B1(_04944_),
    .C1(_04942_),
    .X(_00053_));
 sky130_fd_sc_hd__or2_1 _11877_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][15] ),
    .B(_04943_),
    .X(_04945_));
 sky130_fd_sc_hd__o211a_1 _11878_ (.A1(net544),
    .A2(_04938_),
    .B1(_04945_),
    .C1(_04942_),
    .X(_00054_));
 sky130_fd_sc_hd__or2_1 _11879_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][16] ),
    .B(_04943_),
    .X(_04946_));
 sky130_fd_sc_hd__o211a_1 _11880_ (.A1(net411),
    .A2(_04938_),
    .B1(_04946_),
    .C1(_04942_),
    .X(_00055_));
 sky130_fd_sc_hd__or2_1 _11881_ (.A(net576),
    .B(_04943_),
    .X(_04947_));
 sky130_fd_sc_hd__o211a_1 _11882_ (.A1(net891),
    .A2(_04938_),
    .B1(_04947_),
    .C1(_04942_),
    .X(_00056_));
 sky130_fd_sc_hd__or2_1 _11883_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][18] ),
    .B(_04943_),
    .X(_04948_));
 sky130_fd_sc_hd__o211a_1 _11884_ (.A1(net503),
    .A2(_04938_),
    .B1(_04948_),
    .C1(_04942_),
    .X(_00057_));
 sky130_fd_sc_hd__or2_1 _11885_ (.A(net800),
    .B(_04943_),
    .X(_04949_));
 sky130_fd_sc_hd__o211a_1 _11886_ (.A1(net878),
    .A2(_04938_),
    .B1(_04949_),
    .C1(_04942_),
    .X(_00058_));
 sky130_fd_sc_hd__or2_1 _11887_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][20] ),
    .B(_04943_),
    .X(_04950_));
 sky130_fd_sc_hd__o211a_1 _11888_ (.A1(net886),
    .A2(_04938_),
    .B1(_04950_),
    .C1(_04942_),
    .X(_00059_));
 sky130_fd_sc_hd__clkbuf_4 _11889_ (.A(_04911_),
    .X(_04951_));
 sky130_fd_sc_hd__or2_1 _11890_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][21] ),
    .B(_04943_),
    .X(_04952_));
 sky130_fd_sc_hd__o211a_1 _11891_ (.A1(net648),
    .A2(_04951_),
    .B1(_04952_),
    .C1(_04942_),
    .X(_00060_));
 sky130_fd_sc_hd__or2_1 _11892_ (.A(net474),
    .B(_04943_),
    .X(_04953_));
 sky130_fd_sc_hd__o211a_1 _11893_ (.A1(net636),
    .A2(_04951_),
    .B1(_04953_),
    .C1(_04942_),
    .X(_00061_));
 sky130_fd_sc_hd__or2_1 _11894_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][23] ),
    .B(_04943_),
    .X(_04954_));
 sky130_fd_sc_hd__clkbuf_4 _11895_ (.A(_04874_),
    .X(_04955_));
 sky130_fd_sc_hd__o211a_1 _11896_ (.A1(net670),
    .A2(_04951_),
    .B1(_04954_),
    .C1(_04955_),
    .X(_00062_));
 sky130_fd_sc_hd__clkbuf_4 _11897_ (.A(_04876_),
    .X(_04956_));
 sky130_fd_sc_hd__or2_1 _11898_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][24] ),
    .B(_04956_),
    .X(_04957_));
 sky130_fd_sc_hd__o211a_1 _11899_ (.A1(net524),
    .A2(_04951_),
    .B1(_04957_),
    .C1(_04955_),
    .X(_00063_));
 sky130_fd_sc_hd__or2_1 _11900_ (.A(net652),
    .B(_04956_),
    .X(_04958_));
 sky130_fd_sc_hd__o211a_1 _11901_ (.A1(net953),
    .A2(_04951_),
    .B1(_04958_),
    .C1(_04955_),
    .X(_00064_));
 sky130_fd_sc_hd__or2_1 _11902_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][26] ),
    .B(_04956_),
    .X(_04959_));
 sky130_fd_sc_hd__o211a_1 _11903_ (.A1(net430),
    .A2(_04951_),
    .B1(_04959_),
    .C1(_04955_),
    .X(_00065_));
 sky130_fd_sc_hd__or2_1 _11904_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][27] ),
    .B(_04956_),
    .X(_04960_));
 sky130_fd_sc_hd__o211a_1 _11905_ (.A1(net682),
    .A2(_04951_),
    .B1(_04960_),
    .C1(_04955_),
    .X(_00066_));
 sky130_fd_sc_hd__or2_1 _11906_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][28] ),
    .B(_04956_),
    .X(_04961_));
 sky130_fd_sc_hd__o211a_1 _11907_ (.A1(net668),
    .A2(_04951_),
    .B1(_04961_),
    .C1(_04955_),
    .X(_00067_));
 sky130_fd_sc_hd__or2_1 _11908_ (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][29] ),
    .B(_04956_),
    .X(_04962_));
 sky130_fd_sc_hd__o211a_1 _11909_ (.A1(net561),
    .A2(_04951_),
    .B1(_04962_),
    .C1(_04955_),
    .X(_00068_));
 sky130_fd_sc_hd__or2_1 _11910_ (.A(net689),
    .B(_04956_),
    .X(_04963_));
 sky130_fd_sc_hd__o211a_1 _11911_ (.A1(net868),
    .A2(_04951_),
    .B1(_04963_),
    .C1(_04955_),
    .X(_00069_));
 sky130_fd_sc_hd__clkbuf_4 _11912_ (.A(_04911_),
    .X(_04964_));
 sky130_fd_sc_hd__or2_1 _11913_ (.A(net428),
    .B(_04956_),
    .X(_04965_));
 sky130_fd_sc_hd__o211a_1 _11914_ (.A1(net954),
    .A2(_04964_),
    .B1(_04965_),
    .C1(_04955_),
    .X(_00070_));
 sky130_fd_sc_hd__or2_1 _11915_ (.A(net493),
    .B(_04956_),
    .X(_04966_));
 sky130_fd_sc_hd__o211a_1 _11916_ (.A1(net717),
    .A2(_04964_),
    .B1(_04966_),
    .C1(_04955_),
    .X(_00071_));
 sky130_fd_sc_hd__or2_1 _11917_ (.A(net673),
    .B(_04956_),
    .X(_04967_));
 sky130_fd_sc_hd__clkbuf_4 _11918_ (.A(_04874_),
    .X(_04968_));
 sky130_fd_sc_hd__o211a_1 _11919_ (.A1(net1001),
    .A2(_04964_),
    .B1(_04967_),
    .C1(_04968_),
    .X(_00072_));
 sky130_fd_sc_hd__buf_2 _11920_ (.A(_04876_),
    .X(_04969_));
 sky130_fd_sc_hd__or2_1 _11921_ (.A(\top_inst.axis_out_inst.out_buff_data[34] ),
    .B(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__o211a_1 _11922_ (.A1(net481),
    .A2(_04964_),
    .B1(_04970_),
    .C1(_04968_),
    .X(_00073_));
 sky130_fd_sc_hd__or2_1 _11923_ (.A(\top_inst.axis_out_inst.out_buff_data[35] ),
    .B(_04969_),
    .X(_04971_));
 sky130_fd_sc_hd__o211a_1 _11924_ (.A1(net478),
    .A2(_04964_),
    .B1(_04971_),
    .C1(_04968_),
    .X(_00074_));
 sky130_fd_sc_hd__or2_1 _11925_ (.A(net378),
    .B(_04969_),
    .X(_04972_));
 sky130_fd_sc_hd__o211a_1 _11926_ (.A1(net558),
    .A2(_04964_),
    .B1(_04972_),
    .C1(_04968_),
    .X(_00075_));
 sky130_fd_sc_hd__or2_1 _11927_ (.A(net676),
    .B(_04969_),
    .X(_04973_));
 sky130_fd_sc_hd__o211a_1 _11928_ (.A1(net892),
    .A2(_04964_),
    .B1(_04973_),
    .C1(_04968_),
    .X(_00076_));
 sky130_fd_sc_hd__or2_1 _11929_ (.A(net845),
    .B(_04969_),
    .X(_04974_));
 sky130_fd_sc_hd__o211a_1 _11930_ (.A1(net970),
    .A2(_04964_),
    .B1(_04974_),
    .C1(_04968_),
    .X(_00077_));
 sky130_fd_sc_hd__or2_1 _11931_ (.A(net665),
    .B(_04969_),
    .X(_04975_));
 sky130_fd_sc_hd__o211a_1 _11932_ (.A1(net880),
    .A2(_04964_),
    .B1(_04975_),
    .C1(_04968_),
    .X(_00078_));
 sky130_fd_sc_hd__or2_1 _11933_ (.A(net595),
    .B(_04969_),
    .X(_04976_));
 sky130_fd_sc_hd__o211a_1 _11934_ (.A1(net905),
    .A2(_04964_),
    .B1(_04976_),
    .C1(_04968_),
    .X(_00079_));
 sky130_fd_sc_hd__clkbuf_4 _11935_ (.A(_04911_),
    .X(_04977_));
 sky130_fd_sc_hd__or2_1 _11936_ (.A(\top_inst.axis_out_inst.out_buff_data[41] ),
    .B(_04969_),
    .X(_04978_));
 sky130_fd_sc_hd__o211a_1 _11937_ (.A1(net520),
    .A2(_04977_),
    .B1(_04978_),
    .C1(_04968_),
    .X(_00080_));
 sky130_fd_sc_hd__or2_1 _11938_ (.A(net613),
    .B(_04969_),
    .X(_04979_));
 sky130_fd_sc_hd__o211a_1 _11939_ (.A1(net999),
    .A2(_04977_),
    .B1(_04979_),
    .C1(_04968_),
    .X(_00081_));
 sky130_fd_sc_hd__or2_1 _11940_ (.A(net610),
    .B(_04969_),
    .X(_04980_));
 sky130_fd_sc_hd__clkbuf_4 _11941_ (.A(_04874_),
    .X(_04981_));
 sky130_fd_sc_hd__o211a_1 _11942_ (.A1(net1012),
    .A2(_04977_),
    .B1(_04980_),
    .C1(_04981_),
    .X(_00082_));
 sky130_fd_sc_hd__buf_2 _11943_ (.A(_04876_),
    .X(_04982_));
 sky130_fd_sc_hd__or2_1 _11944_ (.A(net513),
    .B(_04982_),
    .X(_04983_));
 sky130_fd_sc_hd__o211a_1 _11945_ (.A1(net1021),
    .A2(_04977_),
    .B1(_04983_),
    .C1(_04981_),
    .X(_00083_));
 sky130_fd_sc_hd__or2_1 _11946_ (.A(\top_inst.axis_out_inst.out_buff_data[45] ),
    .B(_04982_),
    .X(_04984_));
 sky130_fd_sc_hd__o211a_1 _11947_ (.A1(net549),
    .A2(_04977_),
    .B1(_04984_),
    .C1(_04981_),
    .X(_00084_));
 sky130_fd_sc_hd__or2_1 _11948_ (.A(net731),
    .B(_04982_),
    .X(_04985_));
 sky130_fd_sc_hd__o211a_1 _11949_ (.A1(net913),
    .A2(_04977_),
    .B1(_04985_),
    .C1(_04981_),
    .X(_00085_));
 sky130_fd_sc_hd__or2_1 _11950_ (.A(net651),
    .B(_04982_),
    .X(_04986_));
 sky130_fd_sc_hd__o211a_1 _11951_ (.A1(net733),
    .A2(_04977_),
    .B1(_04986_),
    .C1(_04981_),
    .X(_00086_));
 sky130_fd_sc_hd__or2_1 _11952_ (.A(net553),
    .B(_04982_),
    .X(_04987_));
 sky130_fd_sc_hd__o211a_1 _11953_ (.A1(net967),
    .A2(_04977_),
    .B1(_04987_),
    .C1(_04981_),
    .X(_00087_));
 sky130_fd_sc_hd__or2_1 _11954_ (.A(net699),
    .B(_04982_),
    .X(_04988_));
 sky130_fd_sc_hd__o211a_1 _11955_ (.A1(net876),
    .A2(_04977_),
    .B1(_04988_),
    .C1(_04981_),
    .X(_00088_));
 sky130_fd_sc_hd__or2_1 _11956_ (.A(net796),
    .B(_04982_),
    .X(_04989_));
 sky130_fd_sc_hd__o211a_1 _11957_ (.A1(net864),
    .A2(_04977_),
    .B1(_04989_),
    .C1(_04981_),
    .X(_00089_));
 sky130_fd_sc_hd__clkbuf_4 _11958_ (.A(_04911_),
    .X(_04990_));
 sky130_fd_sc_hd__or2_1 _11959_ (.A(net693),
    .B(_04982_),
    .X(_04991_));
 sky130_fd_sc_hd__o211a_1 _11960_ (.A1(net783),
    .A2(_04990_),
    .B1(_04991_),
    .C1(_04981_),
    .X(_00090_));
 sky130_fd_sc_hd__or2_1 _11961_ (.A(\top_inst.axis_out_inst.out_buff_data[52] ),
    .B(_04982_),
    .X(_04992_));
 sky130_fd_sc_hd__o211a_1 _11962_ (.A1(net914),
    .A2(_04990_),
    .B1(_04992_),
    .C1(_04981_),
    .X(_00091_));
 sky130_fd_sc_hd__or2_1 _11963_ (.A(\top_inst.axis_out_inst.out_buff_data[53] ),
    .B(_04982_),
    .X(_04993_));
 sky130_fd_sc_hd__clkbuf_4 _11964_ (.A(_04873_),
    .X(_04994_));
 sky130_fd_sc_hd__clkbuf_4 _11965_ (.A(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__o211a_1 _11966_ (.A1(net805),
    .A2(_04990_),
    .B1(_04993_),
    .C1(_04995_),
    .X(_00092_));
 sky130_fd_sc_hd__buf_2 _11967_ (.A(_04876_),
    .X(_04996_));
 sky130_fd_sc_hd__or2_1 _11968_ (.A(net802),
    .B(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__o211a_1 _11969_ (.A1(net849),
    .A2(_04990_),
    .B1(_04997_),
    .C1(_04995_),
    .X(_00093_));
 sky130_fd_sc_hd__or2_1 _11970_ (.A(\top_inst.axis_out_inst.out_buff_data[55] ),
    .B(_04996_),
    .X(_04998_));
 sky130_fd_sc_hd__o211a_1 _11971_ (.A1(net700),
    .A2(_04990_),
    .B1(_04998_),
    .C1(_04995_),
    .X(_00094_));
 sky130_fd_sc_hd__or2_1 _11972_ (.A(\top_inst.axis_out_inst.out_buff_data[56] ),
    .B(_04996_),
    .X(_04999_));
 sky130_fd_sc_hd__o211a_1 _11973_ (.A1(net814),
    .A2(_04990_),
    .B1(_04999_),
    .C1(_04995_),
    .X(_00095_));
 sky130_fd_sc_hd__or2_1 _11974_ (.A(\top_inst.axis_out_inst.out_buff_data[57] ),
    .B(_04996_),
    .X(_05000_));
 sky130_fd_sc_hd__o211a_1 _11975_ (.A1(net791),
    .A2(_04990_),
    .B1(_05000_),
    .C1(_04995_),
    .X(_00096_));
 sky130_fd_sc_hd__or2_1 _11976_ (.A(net1101),
    .B(_04996_),
    .X(_05001_));
 sky130_fd_sc_hd__o211a_1 _11977_ (.A1(net973),
    .A2(_04990_),
    .B1(_05001_),
    .C1(_04995_),
    .X(_00097_));
 sky130_fd_sc_hd__or2_1 _11978_ (.A(\top_inst.axis_out_inst.out_buff_data[59] ),
    .B(_04996_),
    .X(_05002_));
 sky130_fd_sc_hd__o211a_1 _11979_ (.A1(net720),
    .A2(_04990_),
    .B1(_05002_),
    .C1(_04995_),
    .X(_00098_));
 sky130_fd_sc_hd__or2_1 _11980_ (.A(\top_inst.axis_out_inst.out_buff_data[60] ),
    .B(_04996_),
    .X(_05003_));
 sky130_fd_sc_hd__o211a_1 _11981_ (.A1(net551),
    .A2(_04990_),
    .B1(_05003_),
    .C1(_04995_),
    .X(_00099_));
 sky130_fd_sc_hd__clkbuf_4 _11982_ (.A(_04911_),
    .X(_05004_));
 sky130_fd_sc_hd__or2_1 _11983_ (.A(\top_inst.axis_out_inst.out_buff_data[61] ),
    .B(_04996_),
    .X(_05005_));
 sky130_fd_sc_hd__o211a_1 _11984_ (.A1(net598),
    .A2(_05004_),
    .B1(_05005_),
    .C1(_04995_),
    .X(_00100_));
 sky130_fd_sc_hd__or2_1 _11985_ (.A(net730),
    .B(_04996_),
    .X(_05006_));
 sky130_fd_sc_hd__o211a_1 _11986_ (.A1(net820),
    .A2(_05004_),
    .B1(_05006_),
    .C1(_04995_),
    .X(_00101_));
 sky130_fd_sc_hd__or2_1 _11987_ (.A(net1108),
    .B(_04996_),
    .X(_05007_));
 sky130_fd_sc_hd__clkbuf_4 _11988_ (.A(_04994_),
    .X(_05008_));
 sky130_fd_sc_hd__o211a_1 _11989_ (.A1(net722),
    .A2(_05004_),
    .B1(_05007_),
    .C1(_05008_),
    .X(_00102_));
 sky130_fd_sc_hd__clkbuf_4 _11990_ (.A(_04863_),
    .X(_05009_));
 sky130_fd_sc_hd__clkbuf_2 _11991_ (.A(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__or2_1 _11992_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][0] ),
    .B(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__o211a_1 _11993_ (.A1(net737),
    .A2(_05004_),
    .B1(_05011_),
    .C1(_05008_),
    .X(_00103_));
 sky130_fd_sc_hd__or2_1 _11994_ (.A(net447),
    .B(_05010_),
    .X(_05012_));
 sky130_fd_sc_hd__o211a_1 _11995_ (.A1(net760),
    .A2(_05004_),
    .B1(_05012_),
    .C1(_05008_),
    .X(_00104_));
 sky130_fd_sc_hd__or2_1 _11996_ (.A(net556),
    .B(_05010_),
    .X(_05013_));
 sky130_fd_sc_hd__o211a_1 _11997_ (.A1(net779),
    .A2(_05004_),
    .B1(_05013_),
    .C1(_05008_),
    .X(_00105_));
 sky130_fd_sc_hd__or2_1 _11998_ (.A(net514),
    .B(_05010_),
    .X(_05014_));
 sky130_fd_sc_hd__o211a_1 _11999_ (.A1(net758),
    .A2(_05004_),
    .B1(_05014_),
    .C1(_05008_),
    .X(_00106_));
 sky130_fd_sc_hd__or2_1 _12000_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][4] ),
    .B(_05010_),
    .X(_05015_));
 sky130_fd_sc_hd__o211a_1 _12001_ (.A1(net497),
    .A2(_05004_),
    .B1(_05015_),
    .C1(_05008_),
    .X(_00107_));
 sky130_fd_sc_hd__or2_1 _12002_ (.A(net797),
    .B(_05010_),
    .X(_05016_));
 sky130_fd_sc_hd__o211a_1 _12003_ (.A1(net894),
    .A2(_05004_),
    .B1(_05016_),
    .C1(_05008_),
    .X(_00108_));
 sky130_fd_sc_hd__or2_1 _12004_ (.A(net458),
    .B(_05010_),
    .X(_05017_));
 sky130_fd_sc_hd__o211a_1 _12005_ (.A1(net862),
    .A2(_05004_),
    .B1(_05017_),
    .C1(_05008_),
    .X(_00109_));
 sky130_fd_sc_hd__buf_2 _12006_ (.A(_04911_),
    .X(_05018_));
 sky130_fd_sc_hd__or2_1 _12007_ (.A(net546),
    .B(_05010_),
    .X(_05019_));
 sky130_fd_sc_hd__o211a_1 _12008_ (.A1(net745),
    .A2(_05018_),
    .B1(_05019_),
    .C1(_05008_),
    .X(_00110_));
 sky130_fd_sc_hd__or2_1 _12009_ (.A(net445),
    .B(_05010_),
    .X(_05020_));
 sky130_fd_sc_hd__o211a_1 _12010_ (.A1(net871),
    .A2(_05018_),
    .B1(_05020_),
    .C1(_05008_),
    .X(_00111_));
 sky130_fd_sc_hd__or2_1 _12011_ (.A(net577),
    .B(_05010_),
    .X(_05021_));
 sky130_fd_sc_hd__buf_2 _12012_ (.A(_04994_),
    .X(_05022_));
 sky130_fd_sc_hd__o211a_1 _12013_ (.A1(net883),
    .A2(_05018_),
    .B1(_05021_),
    .C1(_05022_),
    .X(_00112_));
 sky130_fd_sc_hd__clkbuf_2 _12014_ (.A(_05009_),
    .X(_05023_));
 sky130_fd_sc_hd__or2_1 _12015_ (.A(net488),
    .B(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__o211a_1 _12016_ (.A1(net631),
    .A2(_05018_),
    .B1(_05024_),
    .C1(_05022_),
    .X(_00113_));
 sky130_fd_sc_hd__or2_1 _12017_ (.A(net563),
    .B(_05023_),
    .X(_05025_));
 sky130_fd_sc_hd__o211a_1 _12018_ (.A1(net795),
    .A2(_05018_),
    .B1(_05025_),
    .C1(_05022_),
    .X(_00114_));
 sky130_fd_sc_hd__or2_1 _12019_ (.A(net439),
    .B(_05023_),
    .X(_05026_));
 sky130_fd_sc_hd__o211a_1 _12020_ (.A1(net816),
    .A2(_05018_),
    .B1(_05026_),
    .C1(_05022_),
    .X(_00115_));
 sky130_fd_sc_hd__or2_1 _12021_ (.A(net272),
    .B(_05023_),
    .X(_05027_));
 sky130_fd_sc_hd__o211a_1 _12022_ (.A1(net837),
    .A2(_05018_),
    .B1(_05027_),
    .C1(_05022_),
    .X(_00116_));
 sky130_fd_sc_hd__or2_1 _12023_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][14] ),
    .B(_05023_),
    .X(_05028_));
 sky130_fd_sc_hd__o211a_1 _12024_ (.A1(net315),
    .A2(_05018_),
    .B1(_05028_),
    .C1(_05022_),
    .X(_00117_));
 sky130_fd_sc_hd__or2_1 _12025_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][15] ),
    .B(_05023_),
    .X(_05029_));
 sky130_fd_sc_hd__o211a_1 _12026_ (.A1(net278),
    .A2(_05018_),
    .B1(_05029_),
    .C1(_05022_),
    .X(_00118_));
 sky130_fd_sc_hd__or2_1 _12027_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][16] ),
    .B(_05023_),
    .X(_05030_));
 sky130_fd_sc_hd__o211a_1 _12028_ (.A1(net270),
    .A2(_05018_),
    .B1(_05030_),
    .C1(_05022_),
    .X(_00119_));
 sky130_fd_sc_hd__clkbuf_4 _12029_ (.A(_04911_),
    .X(_05031_));
 sky130_fd_sc_hd__or2_1 _12030_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][17] ),
    .B(_05023_),
    .X(_05032_));
 sky130_fd_sc_hd__o211a_1 _12031_ (.A1(net280),
    .A2(_05031_),
    .B1(_05032_),
    .C1(_05022_),
    .X(_00120_));
 sky130_fd_sc_hd__or2_1 _12032_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][18] ),
    .B(_05023_),
    .X(_05033_));
 sky130_fd_sc_hd__o211a_1 _12033_ (.A1(net268),
    .A2(_05031_),
    .B1(_05033_),
    .C1(_05022_),
    .X(_00121_));
 sky130_fd_sc_hd__or2_1 _12034_ (.A(net1105),
    .B(_05023_),
    .X(_05034_));
 sky130_fd_sc_hd__buf_2 _12035_ (.A(_04994_),
    .X(_05035_));
 sky130_fd_sc_hd__o211a_1 _12036_ (.A1(net966),
    .A2(_05031_),
    .B1(_05034_),
    .C1(_05035_),
    .X(_00122_));
 sky130_fd_sc_hd__clkbuf_2 _12037_ (.A(_05009_),
    .X(_05036_));
 sky130_fd_sc_hd__or2_1 _12038_ (.A(net262),
    .B(_05036_),
    .X(_05037_));
 sky130_fd_sc_hd__o211a_1 _12039_ (.A1(net861),
    .A2(_05031_),
    .B1(_05037_),
    .C1(_05035_),
    .X(_00123_));
 sky130_fd_sc_hd__or2_1 _12040_ (.A(net469),
    .B(_05036_),
    .X(_05038_));
 sky130_fd_sc_hd__o211a_1 _12041_ (.A1(net782),
    .A2(_05031_),
    .B1(_05038_),
    .C1(_05035_),
    .X(_00124_));
 sky130_fd_sc_hd__or2_1 _12042_ (.A(net510),
    .B(_05036_),
    .X(_05039_));
 sky130_fd_sc_hd__o211a_1 _12043_ (.A1(net672),
    .A2(_05031_),
    .B1(_05039_),
    .C1(_05035_),
    .X(_00125_));
 sky130_fd_sc_hd__or2_1 _12044_ (.A(net264),
    .B(_05036_),
    .X(_05040_));
 sky130_fd_sc_hd__o211a_1 _12045_ (.A1(net647),
    .A2(_05031_),
    .B1(_05040_),
    .C1(_05035_),
    .X(_00126_));
 sky130_fd_sc_hd__or2_1 _12046_ (.A(net385),
    .B(_05036_),
    .X(_05041_));
 sky130_fd_sc_hd__o211a_1 _12047_ (.A1(net696),
    .A2(_05031_),
    .B1(_05041_),
    .C1(_05035_),
    .X(_00127_));
 sky130_fd_sc_hd__or2_1 _12048_ (.A(net793),
    .B(_05036_),
    .X(_05042_));
 sky130_fd_sc_hd__o211a_1 _12049_ (.A1(net919),
    .A2(_05031_),
    .B1(_05042_),
    .C1(_05035_),
    .X(_00128_));
 sky130_fd_sc_hd__or2_1 _12050_ (.A(net274),
    .B(_05036_),
    .X(_05043_));
 sky130_fd_sc_hd__o211a_1 _12051_ (.A1(net477),
    .A2(_05031_),
    .B1(_05043_),
    .C1(_05035_),
    .X(_00129_));
 sky130_fd_sc_hd__buf_4 _12052_ (.A(_04858_),
    .X(_05044_));
 sky130_fd_sc_hd__clkbuf_4 _12053_ (.A(_05044_),
    .X(_05045_));
 sky130_fd_sc_hd__or2_1 _12054_ (.A(net256),
    .B(_05036_),
    .X(_05046_));
 sky130_fd_sc_hd__o211a_1 _12055_ (.A1(net997),
    .A2(_05045_),
    .B1(_05046_),
    .C1(_05035_),
    .X(_00130_));
 sky130_fd_sc_hd__or2_1 _12056_ (.A(net266),
    .B(_05036_),
    .X(_05047_));
 sky130_fd_sc_hd__o211a_1 _12057_ (.A1(net869),
    .A2(_05045_),
    .B1(_05047_),
    .C1(_05035_),
    .X(_00131_));
 sky130_fd_sc_hd__or2_1 _12058_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][29] ),
    .B(_05036_),
    .X(_05048_));
 sky130_fd_sc_hd__buf_2 _12059_ (.A(_04994_),
    .X(_05049_));
 sky130_fd_sc_hd__o211a_1 _12060_ (.A1(net327),
    .A2(_05045_),
    .B1(_05048_),
    .C1(_05049_),
    .X(_00132_));
 sky130_fd_sc_hd__clkbuf_2 _12061_ (.A(_05009_),
    .X(_05050_));
 sky130_fd_sc_hd__or2_1 _12062_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][30] ),
    .B(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__o211a_1 _12063_ (.A1(net559),
    .A2(_05045_),
    .B1(_05051_),
    .C1(_05049_),
    .X(_00133_));
 sky130_fd_sc_hd__or2_1 _12064_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][31] ),
    .B(_05050_),
    .X(_05052_));
 sky130_fd_sc_hd__o211a_1 _12065_ (.A1(net518),
    .A2(_05045_),
    .B1(_05052_),
    .C1(_05049_),
    .X(_00134_));
 sky130_fd_sc_hd__or2_1 _12066_ (.A(net717),
    .B(_05050_),
    .X(_05053_));
 sky130_fd_sc_hd__o211a_1 _12067_ (.A1(net877),
    .A2(_05045_),
    .B1(_05053_),
    .C1(_05049_),
    .X(_00135_));
 sky130_fd_sc_hd__or2_1 _12068_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][1] ),
    .B(_05050_),
    .X(_05054_));
 sky130_fd_sc_hd__o211a_1 _12069_ (.A1(net447),
    .A2(_05045_),
    .B1(_05054_),
    .C1(_05049_),
    .X(_00136_));
 sky130_fd_sc_hd__or2_1 _12070_ (.A(net481),
    .B(_05050_),
    .X(_05055_));
 sky130_fd_sc_hd__o211a_1 _12071_ (.A1(net556),
    .A2(_05045_),
    .B1(_05055_),
    .C1(_05049_),
    .X(_00137_));
 sky130_fd_sc_hd__or2_1 _12072_ (.A(net478),
    .B(_05050_),
    .X(_05056_));
 sky130_fd_sc_hd__o211a_1 _12073_ (.A1(net514),
    .A2(_05045_),
    .B1(_05056_),
    .C1(_05049_),
    .X(_00138_));
 sky130_fd_sc_hd__or2_1 _12074_ (.A(net558),
    .B(_05050_),
    .X(_05057_));
 sky130_fd_sc_hd__o211a_1 _12075_ (.A1(net780),
    .A2(_05045_),
    .B1(_05057_),
    .C1(_05049_),
    .X(_00139_));
 sky130_fd_sc_hd__buf_2 _12076_ (.A(_05044_),
    .X(_05058_));
 sky130_fd_sc_hd__or2_1 _12077_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][5] ),
    .B(_05050_),
    .X(_05059_));
 sky130_fd_sc_hd__o211a_1 _12078_ (.A1(net797),
    .A2(_05058_),
    .B1(_05059_),
    .C1(_05049_),
    .X(_00140_));
 sky130_fd_sc_hd__or2_1 _12079_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][6] ),
    .B(_05050_),
    .X(_05060_));
 sky130_fd_sc_hd__o211a_1 _12080_ (.A1(net458),
    .A2(_05058_),
    .B1(_05060_),
    .C1(_05049_),
    .X(_00141_));
 sky130_fd_sc_hd__or2_1 _12081_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][7] ),
    .B(_05050_),
    .X(_05061_));
 sky130_fd_sc_hd__buf_2 _12082_ (.A(_04994_),
    .X(_05062_));
 sky130_fd_sc_hd__o211a_1 _12083_ (.A1(net546),
    .A2(_05058_),
    .B1(_05061_),
    .C1(_05062_),
    .X(_00142_));
 sky130_fd_sc_hd__clkbuf_2 _12084_ (.A(_05009_),
    .X(_05063_));
 sky130_fd_sc_hd__or2_1 _12085_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][8] ),
    .B(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__o211a_1 _12086_ (.A1(net445),
    .A2(_05058_),
    .B1(_05064_),
    .C1(_05062_),
    .X(_00143_));
 sky130_fd_sc_hd__or2_1 _12087_ (.A(net520),
    .B(_05063_),
    .X(_05065_));
 sky130_fd_sc_hd__o211a_1 _12088_ (.A1(net577),
    .A2(_05058_),
    .B1(_05065_),
    .C1(_05062_),
    .X(_00144_));
 sky130_fd_sc_hd__or2_1 _12089_ (.A(net1100),
    .B(_05063_),
    .X(_05066_));
 sky130_fd_sc_hd__o211a_1 _12090_ (.A1(net488),
    .A2(_05058_),
    .B1(_05066_),
    .C1(_05062_),
    .X(_00145_));
 sky130_fd_sc_hd__or2_1 _12091_ (.A(net1104),
    .B(_05063_),
    .X(_05067_));
 sky130_fd_sc_hd__o211a_1 _12092_ (.A1(net563),
    .A2(_05058_),
    .B1(_05067_),
    .C1(_05062_),
    .X(_00146_));
 sky130_fd_sc_hd__or2_1 _12093_ (.A(net1106),
    .B(_05063_),
    .X(_05068_));
 sky130_fd_sc_hd__o211a_1 _12094_ (.A1(net439),
    .A2(_05058_),
    .B1(_05068_),
    .C1(_05062_),
    .X(_00147_));
 sky130_fd_sc_hd__or2_1 _12095_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][13] ),
    .B(_05063_),
    .X(_05069_));
 sky130_fd_sc_hd__o211a_1 _12096_ (.A1(net272),
    .A2(_05058_),
    .B1(_05069_),
    .C1(_05062_),
    .X(_00148_));
 sky130_fd_sc_hd__or2_1 _12097_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][14] ),
    .B(_05063_),
    .X(_05070_));
 sky130_fd_sc_hd__o211a_1 _12098_ (.A1(net538),
    .A2(_05058_),
    .B1(_05070_),
    .C1(_05062_),
    .X(_00149_));
 sky130_fd_sc_hd__clkbuf_4 _12099_ (.A(_05044_),
    .X(_05071_));
 sky130_fd_sc_hd__or2_1 _12100_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][15] ),
    .B(_05063_),
    .X(_05072_));
 sky130_fd_sc_hd__o211a_1 _12101_ (.A1(net587),
    .A2(_05071_),
    .B1(_05072_),
    .C1(_05062_),
    .X(_00150_));
 sky130_fd_sc_hd__or2_1 _12102_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][16] ),
    .B(_05063_),
    .X(_05073_));
 sky130_fd_sc_hd__o211a_1 _12103_ (.A1(net573),
    .A2(_05071_),
    .B1(_05073_),
    .C1(_05062_),
    .X(_00151_));
 sky130_fd_sc_hd__or2_1 _12104_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][17] ),
    .B(_05063_),
    .X(_05074_));
 sky130_fd_sc_hd__clkbuf_4 _12105_ (.A(_04994_),
    .X(_05075_));
 sky130_fd_sc_hd__o211a_1 _12106_ (.A1(net501),
    .A2(_05071_),
    .B1(_05074_),
    .C1(_05075_),
    .X(_00152_));
 sky130_fd_sc_hd__buf_2 _12107_ (.A(_05009_),
    .X(_05076_));
 sky130_fd_sc_hd__or2_1 _12108_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][18] ),
    .B(_05076_),
    .X(_05077_));
 sky130_fd_sc_hd__o211a_1 _12109_ (.A1(net486),
    .A2(_05071_),
    .B1(_05077_),
    .C1(_05075_),
    .X(_00153_));
 sky130_fd_sc_hd__or2_1 _12110_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][19] ),
    .B(_05076_),
    .X(_05078_));
 sky130_fd_sc_hd__o211a_1 _12111_ (.A1(net254),
    .A2(_05071_),
    .B1(_05078_),
    .C1(_05075_),
    .X(_00154_));
 sky130_fd_sc_hd__or2_1 _12112_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][20] ),
    .B(_05076_),
    .X(_05079_));
 sky130_fd_sc_hd__o211a_1 _12113_ (.A1(net262),
    .A2(_05071_),
    .B1(_05079_),
    .C1(_05075_),
    .X(_00155_));
 sky130_fd_sc_hd__or2_1 _12114_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][21] ),
    .B(_05076_),
    .X(_05080_));
 sky130_fd_sc_hd__o211a_1 _12115_ (.A1(net469),
    .A2(_05071_),
    .B1(_05080_),
    .C1(_05075_),
    .X(_00156_));
 sky130_fd_sc_hd__or2_1 _12116_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][22] ),
    .B(_05076_),
    .X(_05081_));
 sky130_fd_sc_hd__o211a_1 _12117_ (.A1(net510),
    .A2(_05071_),
    .B1(_05081_),
    .C1(_05075_),
    .X(_00157_));
 sky130_fd_sc_hd__or2_1 _12118_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][23] ),
    .B(_05076_),
    .X(_05082_));
 sky130_fd_sc_hd__o211a_1 _12119_ (.A1(net264),
    .A2(_05071_),
    .B1(_05082_),
    .C1(_05075_),
    .X(_00158_));
 sky130_fd_sc_hd__or2_1 _12120_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][24] ),
    .B(_05076_),
    .X(_05083_));
 sky130_fd_sc_hd__o211a_1 _12121_ (.A1(net385),
    .A2(_05071_),
    .B1(_05083_),
    .C1(_05075_),
    .X(_00159_));
 sky130_fd_sc_hd__clkbuf_4 _12122_ (.A(_05044_),
    .X(_05084_));
 sky130_fd_sc_hd__or2_1 _12123_ (.A(net791),
    .B(_05076_),
    .X(_05085_));
 sky130_fd_sc_hd__o211a_1 _12124_ (.A1(net793),
    .A2(_05084_),
    .B1(_05085_),
    .C1(_05075_),
    .X(_00160_));
 sky130_fd_sc_hd__or2_1 _12125_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][26] ),
    .B(_05076_),
    .X(_05086_));
 sky130_fd_sc_hd__o211a_1 _12126_ (.A1(net274),
    .A2(_05084_),
    .B1(_05086_),
    .C1(_05075_),
    .X(_00161_));
 sky130_fd_sc_hd__or2_1 _12127_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][27] ),
    .B(_05076_),
    .X(_05087_));
 sky130_fd_sc_hd__clkbuf_4 _12128_ (.A(_04994_),
    .X(_05088_));
 sky130_fd_sc_hd__o211a_1 _12129_ (.A1(net256),
    .A2(_05084_),
    .B1(_05087_),
    .C1(_05088_),
    .X(_00162_));
 sky130_fd_sc_hd__buf_2 _12130_ (.A(_05009_),
    .X(_05089_));
 sky130_fd_sc_hd__or2_1 _12131_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][28] ),
    .B(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__o211a_1 _12132_ (.A1(net266),
    .A2(_05084_),
    .B1(_05090_),
    .C1(_05088_),
    .X(_00163_));
 sky130_fd_sc_hd__or2_1 _12133_ (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][29] ),
    .B(_05089_),
    .X(_05091_));
 sky130_fd_sc_hd__o211a_1 _12134_ (.A1(net506),
    .A2(_05084_),
    .B1(_05091_),
    .C1(_05088_),
    .X(_00164_));
 sky130_fd_sc_hd__or2_1 _12135_ (.A(net820),
    .B(_05089_),
    .X(_05092_));
 sky130_fd_sc_hd__o211a_1 _12136_ (.A1(net823),
    .A2(_05084_),
    .B1(_05092_),
    .C1(_05088_),
    .X(_00165_));
 sky130_fd_sc_hd__or2_1 _12137_ (.A(net722),
    .B(_05089_),
    .X(_05093_));
 sky130_fd_sc_hd__o211a_1 _12138_ (.A1(net854),
    .A2(_05084_),
    .B1(_05093_),
    .C1(_05088_),
    .X(_00166_));
 sky130_fd_sc_hd__or2_1 _12139_ (.A(\top_inst.axis_out_inst.out_buff_data[0] ),
    .B(_05089_),
    .X(_05094_));
 sky130_fd_sc_hd__o211a_1 _12140_ (.A1(net930),
    .A2(_05084_),
    .B1(_05094_),
    .C1(_05088_),
    .X(_00167_));
 sky130_fd_sc_hd__or2_1 _12141_ (.A(\top_inst.axis_out_inst.out_buff_data[1] ),
    .B(_05089_),
    .X(_05095_));
 sky130_fd_sc_hd__o211a_1 _12142_ (.A1(net432),
    .A2(_05084_),
    .B1(_05095_),
    .C1(_05088_),
    .X(_00168_));
 sky130_fd_sc_hd__or2_1 _12143_ (.A(net677),
    .B(_05089_),
    .X(_05096_));
 sky130_fd_sc_hd__o211a_1 _12144_ (.A1(net835),
    .A2(_05084_),
    .B1(_05096_),
    .C1(_05088_),
    .X(_00169_));
 sky130_fd_sc_hd__clkbuf_4 _12145_ (.A(_05044_),
    .X(_05097_));
 sky130_fd_sc_hd__or2_1 _12146_ (.A(net463),
    .B(_05089_),
    .X(_05098_));
 sky130_fd_sc_hd__o211a_1 _12147_ (.A1(net750),
    .A2(_05097_),
    .B1(_05098_),
    .C1(_05088_),
    .X(_00170_));
 sky130_fd_sc_hd__or2_1 _12148_ (.A(\top_inst.axis_out_inst.out_buff_data[4] ),
    .B(_05089_),
    .X(_05099_));
 sky130_fd_sc_hd__o211a_1 _12149_ (.A1(net398),
    .A2(_05097_),
    .B1(_05099_),
    .C1(_05088_),
    .X(_00171_));
 sky130_fd_sc_hd__or2_1 _12150_ (.A(net686),
    .B(_05089_),
    .X(_05100_));
 sky130_fd_sc_hd__clkbuf_4 _12151_ (.A(_04994_),
    .X(_05101_));
 sky130_fd_sc_hd__o211a_1 _12152_ (.A1(net741),
    .A2(_05097_),
    .B1(_05100_),
    .C1(_05101_),
    .X(_00172_));
 sky130_fd_sc_hd__buf_2 _12153_ (.A(_05009_),
    .X(_05102_));
 sky130_fd_sc_hd__or2_1 _12154_ (.A(\top_inst.axis_out_inst.out_buff_data[6] ),
    .B(_05102_),
    .X(_05103_));
 sky130_fd_sc_hd__o211a_1 _12155_ (.A1(net402),
    .A2(_05097_),
    .B1(_05103_),
    .C1(_05101_),
    .X(_00173_));
 sky130_fd_sc_hd__or2_1 _12156_ (.A(\top_inst.axis_out_inst.out_buff_data[7] ),
    .B(_05102_),
    .X(_05104_));
 sky130_fd_sc_hd__o211a_1 _12157_ (.A1(net418),
    .A2(_05097_),
    .B1(_05104_),
    .C1(_05101_),
    .X(_00174_));
 sky130_fd_sc_hd__or2_1 _12158_ (.A(net310),
    .B(_05102_),
    .X(_05105_));
 sky130_fd_sc_hd__o211a_1 _12159_ (.A1(net775),
    .A2(_05097_),
    .B1(_05105_),
    .C1(_05101_),
    .X(_00175_));
 sky130_fd_sc_hd__or2_1 _12160_ (.A(\top_inst.axis_out_inst.out_buff_data[9] ),
    .B(_05102_),
    .X(_05106_));
 sky130_fd_sc_hd__o211a_1 _12161_ (.A1(net373),
    .A2(_05097_),
    .B1(_05106_),
    .C1(_05101_),
    .X(_00176_));
 sky130_fd_sc_hd__or2_1 _12162_ (.A(\top_inst.axis_out_inst.out_buff_data[10] ),
    .B(_05102_),
    .X(_05107_));
 sky130_fd_sc_hd__o211a_1 _12163_ (.A1(net357),
    .A2(_05097_),
    .B1(_05107_),
    .C1(_05101_),
    .X(_00177_));
 sky130_fd_sc_hd__or2_1 _12164_ (.A(\top_inst.axis_out_inst.out_buff_data[11] ),
    .B(_05102_),
    .X(_05108_));
 sky130_fd_sc_hd__o211a_1 _12165_ (.A1(net592),
    .A2(_05097_),
    .B1(_05108_),
    .C1(_05101_),
    .X(_00178_));
 sky130_fd_sc_hd__or2_1 _12166_ (.A(net618),
    .B(_05102_),
    .X(_05109_));
 sky130_fd_sc_hd__o211a_1 _12167_ (.A1(net855),
    .A2(_05097_),
    .B1(_05109_),
    .C1(_05101_),
    .X(_00179_));
 sky130_fd_sc_hd__clkbuf_4 _12168_ (.A(_05044_),
    .X(_05110_));
 sky130_fd_sc_hd__or2_1 _12169_ (.A(net317),
    .B(_05102_),
    .X(_05111_));
 sky130_fd_sc_hd__o211a_1 _12170_ (.A1(net566),
    .A2(_05110_),
    .B1(_05111_),
    .C1(_05101_),
    .X(_00180_));
 sky130_fd_sc_hd__or2_1 _12171_ (.A(net359),
    .B(_05102_),
    .X(_05112_));
 sky130_fd_sc_hd__o211a_1 _12172_ (.A1(net692),
    .A2(_05110_),
    .B1(_05112_),
    .C1(_05101_),
    .X(_00181_));
 sky130_fd_sc_hd__or2_1 _12173_ (.A(\top_inst.axis_out_inst.out_buff_data[15] ),
    .B(_05102_),
    .X(_05113_));
 sky130_fd_sc_hd__clkbuf_4 _12174_ (.A(_04994_),
    .X(_05114_));
 sky130_fd_sc_hd__o211a_1 _12175_ (.A1(net323),
    .A2(_05110_),
    .B1(_05113_),
    .C1(_05114_),
    .X(_00182_));
 sky130_fd_sc_hd__buf_2 _12176_ (.A(_05009_),
    .X(_05115_));
 sky130_fd_sc_hd__or2_1 _12177_ (.A(\top_inst.axis_out_inst.out_buff_data[16] ),
    .B(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__o211a_1 _12178_ (.A1(net346),
    .A2(_05110_),
    .B1(_05116_),
    .C1(_05114_),
    .X(_00183_));
 sky130_fd_sc_hd__or2_1 _12179_ (.A(net485),
    .B(_05115_),
    .X(_05117_));
 sky130_fd_sc_hd__o211a_1 _12180_ (.A1(net885),
    .A2(_05110_),
    .B1(_05117_),
    .C1(_05114_),
    .X(_00184_));
 sky130_fd_sc_hd__or2_1 _12181_ (.A(\top_inst.axis_out_inst.out_buff_data[18] ),
    .B(_05115_),
    .X(_05118_));
 sky130_fd_sc_hd__o211a_1 _12182_ (.A1(net341),
    .A2(_05110_),
    .B1(_05118_),
    .C1(_05114_),
    .X(_00185_));
 sky130_fd_sc_hd__or2_1 _12183_ (.A(\top_inst.axis_out_inst.out_buff_data[19] ),
    .B(_05115_),
    .X(_05119_));
 sky130_fd_sc_hd__o211a_1 _12184_ (.A1(net350),
    .A2(_05110_),
    .B1(_05119_),
    .C1(_05114_),
    .X(_00186_));
 sky130_fd_sc_hd__or2_1 _12185_ (.A(net382),
    .B(_05115_),
    .X(_05120_));
 sky130_fd_sc_hd__o211a_1 _12186_ (.A1(net759),
    .A2(_05110_),
    .B1(_05120_),
    .C1(_05114_),
    .X(_00187_));
 sky130_fd_sc_hd__or2_1 _12187_ (.A(net799),
    .B(_05115_),
    .X(_05121_));
 sky130_fd_sc_hd__o211a_1 _12188_ (.A1(net836),
    .A2(_05110_),
    .B1(_05121_),
    .C1(_05114_),
    .X(_00188_));
 sky130_fd_sc_hd__or2_1 _12189_ (.A(\top_inst.axis_out_inst.out_buff_data[22] ),
    .B(_05115_),
    .X(_05122_));
 sky130_fd_sc_hd__o211a_1 _12190_ (.A1(net352),
    .A2(_05110_),
    .B1(_05122_),
    .C1(_05114_),
    .X(_00189_));
 sky130_fd_sc_hd__clkbuf_4 _12191_ (.A(_05044_),
    .X(_05123_));
 sky130_fd_sc_hd__or2_1 _12192_ (.A(\top_inst.axis_out_inst.out_buff_data[23] ),
    .B(_05115_),
    .X(_05124_));
 sky130_fd_sc_hd__o211a_1 _12193_ (.A1(net365),
    .A2(_05123_),
    .B1(_05124_),
    .C1(_05114_),
    .X(_00190_));
 sky130_fd_sc_hd__or2_1 _12194_ (.A(net379),
    .B(_05115_),
    .X(_05125_));
 sky130_fd_sc_hd__o211a_1 _12195_ (.A1(net900),
    .A2(_05123_),
    .B1(_05125_),
    .C1(_05114_),
    .X(_00191_));
 sky130_fd_sc_hd__or2_1 _12196_ (.A(\top_inst.axis_out_inst.out_buff_data[25] ),
    .B(_05115_),
    .X(_05126_));
 sky130_fd_sc_hd__buf_2 _12197_ (.A(_04873_),
    .X(_05127_));
 sky130_fd_sc_hd__clkbuf_4 _12198_ (.A(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__o211a_1 _12199_ (.A1(net526),
    .A2(_05123_),
    .B1(_05126_),
    .C1(_05128_),
    .X(_00192_));
 sky130_fd_sc_hd__buf_2 _12200_ (.A(_05009_),
    .X(_05129_));
 sky130_fd_sc_hd__or2_1 _12201_ (.A(net723),
    .B(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__o211a_1 _12202_ (.A1(net910),
    .A2(_05123_),
    .B1(_05130_),
    .C1(_05128_),
    .X(_00193_));
 sky130_fd_sc_hd__or2_1 _12203_ (.A(net768),
    .B(_05129_),
    .X(_05131_));
 sky130_fd_sc_hd__o211a_1 _12204_ (.A1(net895),
    .A2(_05123_),
    .B1(_05131_),
    .C1(_05128_),
    .X(_00194_));
 sky130_fd_sc_hd__or2_1 _12205_ (.A(\top_inst.axis_out_inst.out_buff_data[28] ),
    .B(_05129_),
    .X(_05132_));
 sky130_fd_sc_hd__o211a_1 _12206_ (.A1(net308),
    .A2(_05123_),
    .B1(_05132_),
    .C1(_05128_),
    .X(_00195_));
 sky130_fd_sc_hd__or2_1 _12207_ (.A(\top_inst.axis_out_inst.out_buff_data[29] ),
    .B(_05129_),
    .X(_05133_));
 sky130_fd_sc_hd__o211a_1 _12208_ (.A1(net375),
    .A2(_05123_),
    .B1(_05133_),
    .C1(_05128_),
    .X(_00196_));
 sky130_fd_sc_hd__or2_1 _12209_ (.A(\top_inst.axis_out_inst.out_buff_data[30] ),
    .B(_05129_),
    .X(_05134_));
 sky130_fd_sc_hd__o211a_1 _12210_ (.A1(net339),
    .A2(_05123_),
    .B1(_05134_),
    .C1(_05128_),
    .X(_00197_));
 sky130_fd_sc_hd__or2_1 _12211_ (.A(\top_inst.axis_out_inst.out_buff_data[31] ),
    .B(_05129_),
    .X(_05135_));
 sky130_fd_sc_hd__o211a_1 _12212_ (.A1(net383),
    .A2(_05123_),
    .B1(_05135_),
    .C1(_05128_),
    .X(_00198_));
 sky130_fd_sc_hd__or2_1 _12213_ (.A(net589),
    .B(_05129_),
    .X(_05136_));
 sky130_fd_sc_hd__o211a_1 _12214_ (.A1(net917),
    .A2(_05123_),
    .B1(_05136_),
    .C1(_05128_),
    .X(_00199_));
 sky130_fd_sc_hd__clkbuf_4 _12215_ (.A(_05044_),
    .X(_05137_));
 sky130_fd_sc_hd__or2_1 _12216_ (.A(net642),
    .B(_05129_),
    .X(_05138_));
 sky130_fd_sc_hd__o211a_1 _12217_ (.A1(net932),
    .A2(_05137_),
    .B1(_05138_),
    .C1(_05128_),
    .X(_00200_));
 sky130_fd_sc_hd__or2_1 _12218_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][2] ),
    .B(_05129_),
    .X(_05139_));
 sky130_fd_sc_hd__o211a_1 _12219_ (.A1(net408),
    .A2(_05137_),
    .B1(_05139_),
    .C1(_05128_),
    .X(_00201_));
 sky130_fd_sc_hd__or2_1 _12220_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][3] ),
    .B(_05129_),
    .X(_05140_));
 sky130_fd_sc_hd__buf_2 _12221_ (.A(_05127_),
    .X(_05141_));
 sky130_fd_sc_hd__o211a_1 _12222_ (.A1(net343),
    .A2(_05137_),
    .B1(_05140_),
    .C1(_05141_),
    .X(_00202_));
 sky130_fd_sc_hd__clkbuf_4 _12223_ (.A(_04863_),
    .X(_05142_));
 sky130_fd_sc_hd__clkbuf_2 _12224_ (.A(_05142_),
    .X(_05143_));
 sky130_fd_sc_hd__or2_1 _12225_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][4] ),
    .B(_05143_),
    .X(_05144_));
 sky130_fd_sc_hd__o211a_1 _12226_ (.A1(net355),
    .A2(_05137_),
    .B1(_05144_),
    .C1(_05141_),
    .X(_00203_));
 sky130_fd_sc_hd__or2_1 _12227_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][5] ),
    .B(_05143_),
    .X(_05145_));
 sky130_fd_sc_hd__o211a_1 _12228_ (.A1(net812),
    .A2(_05137_),
    .B1(_05145_),
    .C1(_05141_),
    .X(_00204_));
 sky130_fd_sc_hd__or2_1 _12229_ (.A(net554),
    .B(_05143_),
    .X(_05146_));
 sky130_fd_sc_hd__o211a_1 _12230_ (.A1(net911),
    .A2(_05137_),
    .B1(_05146_),
    .C1(_05141_),
    .X(_00205_));
 sky130_fd_sc_hd__or2_1 _12231_ (.A(net528),
    .B(_05143_),
    .X(_05147_));
 sky130_fd_sc_hd__o211a_1 _12232_ (.A1(net585),
    .A2(_05137_),
    .B1(_05147_),
    .C1(_05141_),
    .X(_00206_));
 sky130_fd_sc_hd__or2_1 _12233_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][8] ),
    .B(_05143_),
    .X(_05148_));
 sky130_fd_sc_hd__o211a_1 _12234_ (.A1(net846),
    .A2(_05137_),
    .B1(_05148_),
    .C1(_05141_),
    .X(_00207_));
 sky130_fd_sc_hd__or2_1 _12235_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][9] ),
    .B(_05143_),
    .X(_05149_));
 sky130_fd_sc_hd__o211a_1 _12236_ (.A1(net464),
    .A2(_05137_),
    .B1(_05149_),
    .C1(_05141_),
    .X(_00208_));
 sky130_fd_sc_hd__or2_1 _12237_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][10] ),
    .B(_05143_),
    .X(_05150_));
 sky130_fd_sc_hd__o211a_1 _12238_ (.A1(net426),
    .A2(_05137_),
    .B1(_05150_),
    .C1(_05141_),
    .X(_00209_));
 sky130_fd_sc_hd__clkbuf_4 _12239_ (.A(_05044_),
    .X(_05151_));
 sky130_fd_sc_hd__or2_1 _12240_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][11] ),
    .B(_05143_),
    .X(_05152_));
 sky130_fd_sc_hd__o211a_1 _12241_ (.A1(net420),
    .A2(_05151_),
    .B1(_05152_),
    .C1(_05141_),
    .X(_00210_));
 sky130_fd_sc_hd__or2_1 _12242_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][12] ),
    .B(_05143_),
    .X(_05153_));
 sky130_fd_sc_hd__o211a_1 _12243_ (.A1(net826),
    .A2(_05151_),
    .B1(_05153_),
    .C1(_05141_),
    .X(_00211_));
 sky130_fd_sc_hd__or2_1 _12244_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][13] ),
    .B(_05143_),
    .X(_05154_));
 sky130_fd_sc_hd__buf_2 _12245_ (.A(_05127_),
    .X(_05155_));
 sky130_fd_sc_hd__o211a_1 _12246_ (.A1(net596),
    .A2(_05151_),
    .B1(_05154_),
    .C1(_05155_),
    .X(_00212_));
 sky130_fd_sc_hd__clkbuf_2 _12247_ (.A(_05142_),
    .X(_05156_));
 sky130_fd_sc_hd__or2_1 _12248_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][14] ),
    .B(_05156_),
    .X(_05157_));
 sky130_fd_sc_hd__o211a_1 _12249_ (.A1(net483),
    .A2(_05151_),
    .B1(_05157_),
    .C1(_05155_),
    .X(_00213_));
 sky130_fd_sc_hd__or2_1 _12250_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][15] ),
    .B(_05156_),
    .X(_05158_));
 sky130_fd_sc_hd__o211a_1 _12251_ (.A1(net437),
    .A2(_05151_),
    .B1(_05158_),
    .C1(_05155_),
    .X(_00214_));
 sky130_fd_sc_hd__or2_1 _12252_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][16] ),
    .B(_05156_),
    .X(_05159_));
 sky130_fd_sc_hd__o211a_1 _12253_ (.A1(net311),
    .A2(_05151_),
    .B1(_05159_),
    .C1(_05155_),
    .X(_00215_));
 sky130_fd_sc_hd__or2_1 _12254_ (.A(net586),
    .B(_05156_),
    .X(_05160_));
 sky130_fd_sc_hd__o211a_1 _12255_ (.A1(net968),
    .A2(_05151_),
    .B1(_05160_),
    .C1(_05155_),
    .X(_00216_));
 sky130_fd_sc_hd__or2_1 _12256_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][18] ),
    .B(_05156_),
    .X(_05161_));
 sky130_fd_sc_hd__o211a_1 _12257_ (.A1(net435),
    .A2(_05151_),
    .B1(_05161_),
    .C1(_05155_),
    .X(_00217_));
 sky130_fd_sc_hd__or2_1 _12258_ (.A(net863),
    .B(_05156_),
    .X(_05162_));
 sky130_fd_sc_hd__o211a_1 _12259_ (.A1(net907),
    .A2(_05151_),
    .B1(_05162_),
    .C1(_05155_),
    .X(_00218_));
 sky130_fd_sc_hd__or2_1 _12260_ (.A(net678),
    .B(_05156_),
    .X(_05163_));
 sky130_fd_sc_hd__o211a_1 _12261_ (.A1(net925),
    .A2(_05151_),
    .B1(_05163_),
    .C1(_05155_),
    .X(_00219_));
 sky130_fd_sc_hd__buf_2 _12262_ (.A(_05044_),
    .X(_05164_));
 sky130_fd_sc_hd__or2_1 _12263_ (.A(net540),
    .B(_05156_),
    .X(_05165_));
 sky130_fd_sc_hd__o211a_1 _12264_ (.A1(net958),
    .A2(_05164_),
    .B1(_05165_),
    .C1(_05155_),
    .X(_00220_));
 sky130_fd_sc_hd__or2_1 _12265_ (.A(net650),
    .B(_05156_),
    .X(_05166_));
 sky130_fd_sc_hd__o211a_1 _12266_ (.A1(net825),
    .A2(_05164_),
    .B1(_05166_),
    .C1(_05155_),
    .X(_00221_));
 sky130_fd_sc_hd__or2_1 _12267_ (.A(net726),
    .B(_05156_),
    .X(_05167_));
 sky130_fd_sc_hd__buf_2 _12268_ (.A(_05127_),
    .X(_05168_));
 sky130_fd_sc_hd__o211a_1 _12269_ (.A1(net934),
    .A2(_05164_),
    .B1(_05167_),
    .C1(_05168_),
    .X(_00222_));
 sky130_fd_sc_hd__buf_2 _12270_ (.A(_05142_),
    .X(_05169_));
 sky130_fd_sc_hd__or2_1 _12271_ (.A(net698),
    .B(_05169_),
    .X(_05170_));
 sky130_fd_sc_hd__o211a_1 _12272_ (.A1(net786),
    .A2(_05164_),
    .B1(_05170_),
    .C1(_05168_),
    .X(_00223_));
 sky130_fd_sc_hd__or2_1 _12273_ (.A(net879),
    .B(_05169_),
    .X(_05171_));
 sky130_fd_sc_hd__o211a_1 _12274_ (.A1(net976),
    .A2(_05164_),
    .B1(_05171_),
    .C1(_05168_),
    .X(_00224_));
 sky130_fd_sc_hd__or2_1 _12275_ (.A(net747),
    .B(_05169_),
    .X(_05172_));
 sky130_fd_sc_hd__o211a_1 _12276_ (.A1(net906),
    .A2(_05164_),
    .B1(_05172_),
    .C1(_05168_),
    .X(_00225_));
 sky130_fd_sc_hd__or2_1 _12277_ (.A(net306),
    .B(_05169_),
    .X(_05173_));
 sky130_fd_sc_hd__o211a_1 _12278_ (.A1(net981),
    .A2(_05164_),
    .B1(_05173_),
    .C1(_05168_),
    .X(_00226_));
 sky130_fd_sc_hd__or2_1 _12279_ (.A(net691),
    .B(_05169_),
    .X(_05174_));
 sky130_fd_sc_hd__o211a_1 _12280_ (.A1(net756),
    .A2(_05164_),
    .B1(_05174_),
    .C1(_05168_),
    .X(_00227_));
 sky130_fd_sc_hd__or2_1 _12281_ (.A(net695),
    .B(_05169_),
    .X(_05175_));
 sky130_fd_sc_hd__o211a_1 _12282_ (.A1(net790),
    .A2(_05164_),
    .B1(_05175_),
    .C1(_05168_),
    .X(_00228_));
 sky130_fd_sc_hd__or2_1 _12283_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][30] ),
    .B(_05169_),
    .X(_05176_));
 sky130_fd_sc_hd__o211a_1 _12284_ (.A1(net400),
    .A2(_05164_),
    .B1(_05176_),
    .C1(_05168_),
    .X(_00229_));
 sky130_fd_sc_hd__clkbuf_8 _12285_ (.A(_04858_),
    .X(_05177_));
 sky130_fd_sc_hd__clkbuf_4 _12286_ (.A(_05177_),
    .X(_05178_));
 sky130_fd_sc_hd__or2_1 _12287_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][31] ),
    .B(_05169_),
    .X(_05179_));
 sky130_fd_sc_hd__o211a_1 _12288_ (.A1(net490),
    .A2(_05178_),
    .B1(_05179_),
    .C1(_05168_),
    .X(_00230_));
 sky130_fd_sc_hd__or2_1 _12289_ (.A(net495),
    .B(_05169_),
    .X(_05180_));
 sky130_fd_sc_hd__o211a_1 _12290_ (.A1(net589),
    .A2(_05178_),
    .B1(_05180_),
    .C1(_05168_),
    .X(_00231_));
 sky130_fd_sc_hd__or2_1 _12291_ (.A(net466),
    .B(_05169_),
    .X(_05181_));
 sky130_fd_sc_hd__buf_2 _12292_ (.A(_05127_),
    .X(_05182_));
 sky130_fd_sc_hd__o211a_1 _12293_ (.A1(net642),
    .A2(_05178_),
    .B1(_05181_),
    .C1(_05182_),
    .X(_00232_));
 sky130_fd_sc_hd__clkbuf_2 _12294_ (.A(_05142_),
    .X(_05183_));
 sky130_fd_sc_hd__or2_1 _12295_ (.A(net848),
    .B(_05183_),
    .X(_05184_));
 sky130_fd_sc_hd__o211a_1 _12296_ (.A1(net858),
    .A2(_05178_),
    .B1(_05184_),
    .C1(_05182_),
    .X(_00233_));
 sky130_fd_sc_hd__or2_1 _12297_ (.A(net456),
    .B(_05183_),
    .X(_05185_));
 sky130_fd_sc_hd__o211a_1 _12298_ (.A1(net494),
    .A2(_05178_),
    .B1(_05185_),
    .C1(_05182_),
    .X(_00234_));
 sky130_fd_sc_hd__or2_1 _12299_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][4] ),
    .B(_05183_),
    .X(_05186_));
 sky130_fd_sc_hd__o211a_1 _12300_ (.A1(net600),
    .A2(_05178_),
    .B1(_05186_),
    .C1(_05182_),
    .X(_00235_));
 sky130_fd_sc_hd__or2_1 _12301_ (.A(net452),
    .B(_05183_),
    .X(_05187_));
 sky130_fd_sc_hd__o211a_1 _12302_ (.A1(net874),
    .A2(_05178_),
    .B1(_05187_),
    .C1(_05182_),
    .X(_00236_));
 sky130_fd_sc_hd__or2_1 _12303_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][6] ),
    .B(_05183_),
    .X(_05188_));
 sky130_fd_sc_hd__o211a_1 _12304_ (.A1(net554),
    .A2(_05178_),
    .B1(_05188_),
    .C1(_05182_),
    .X(_00237_));
 sky130_fd_sc_hd__or2_1 _12305_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][7] ),
    .B(_05183_),
    .X(_05189_));
 sky130_fd_sc_hd__o211a_1 _12306_ (.A1(net528),
    .A2(_05178_),
    .B1(_05189_),
    .C1(_05182_),
    .X(_00238_));
 sky130_fd_sc_hd__or2_1 _12307_ (.A(net568),
    .B(_05183_),
    .X(_05190_));
 sky130_fd_sc_hd__o211a_1 _12308_ (.A1(net909),
    .A2(_05178_),
    .B1(_05190_),
    .C1(_05182_),
    .X(_00239_));
 sky130_fd_sc_hd__buf_2 _12309_ (.A(_05177_),
    .X(_05191_));
 sky130_fd_sc_hd__or2_1 _12310_ (.A(net572),
    .B(_05183_),
    .X(_05192_));
 sky130_fd_sc_hd__o211a_1 _12311_ (.A1(net916),
    .A2(_05191_),
    .B1(_05192_),
    .C1(_05182_),
    .X(_00240_));
 sky130_fd_sc_hd__or2_1 _12312_ (.A(net807),
    .B(_05183_),
    .X(_05193_));
 sky130_fd_sc_hd__o211a_1 _12313_ (.A1(net841),
    .A2(_05191_),
    .B1(_05193_),
    .C1(_05182_),
    .X(_00241_));
 sky130_fd_sc_hd__or2_1 _12314_ (.A(net535),
    .B(_05183_),
    .X(_05194_));
 sky130_fd_sc_hd__buf_2 _12315_ (.A(_05127_),
    .X(_05195_));
 sky130_fd_sc_hd__o211a_1 _12316_ (.A1(net875),
    .A2(_05191_),
    .B1(_05194_),
    .C1(_05195_),
    .X(_00242_));
 sky130_fd_sc_hd__clkbuf_2 _12317_ (.A(_05142_),
    .X(_05196_));
 sky130_fd_sc_hd__or2_1 _12318_ (.A(net449),
    .B(_05196_),
    .X(_05197_));
 sky130_fd_sc_hd__o211a_1 _12319_ (.A1(net941),
    .A2(_05191_),
    .B1(_05197_),
    .C1(_05195_),
    .X(_00243_));
 sky130_fd_sc_hd__or2_1 _12320_ (.A(net567),
    .B(_05196_),
    .X(_05198_));
 sky130_fd_sc_hd__o211a_1 _12321_ (.A1(net824),
    .A2(_05191_),
    .B1(_05198_),
    .C1(_05195_),
    .X(_00244_));
 sky130_fd_sc_hd__or2_1 _12322_ (.A(net515),
    .B(_05196_),
    .X(_05199_));
 sky130_fd_sc_hd__o211a_1 _12323_ (.A1(net926),
    .A2(_05191_),
    .B1(_05199_),
    .C1(_05195_),
    .X(_00245_));
 sky130_fd_sc_hd__or2_1 _12324_ (.A(net505),
    .B(_05196_),
    .X(_05200_));
 sky130_fd_sc_hd__o211a_1 _12325_ (.A1(net943),
    .A2(_05191_),
    .B1(_05200_),
    .C1(_05195_),
    .X(_00246_));
 sky130_fd_sc_hd__or2_1 _12326_ (.A(net480),
    .B(_05196_),
    .X(_05201_));
 sky130_fd_sc_hd__o211a_1 _12327_ (.A1(net890),
    .A2(_05191_),
    .B1(_05201_),
    .C1(_05195_),
    .X(_00247_));
 sky130_fd_sc_hd__or2_1 _12328_ (.A(net319),
    .B(_05196_),
    .X(_05202_));
 sky130_fd_sc_hd__o211a_1 _12329_ (.A1(net586),
    .A2(_05191_),
    .B1(_05202_),
    .C1(_05195_),
    .X(_00248_));
 sky130_fd_sc_hd__or2_1 _12330_ (.A(net345),
    .B(_05196_),
    .X(_05203_));
 sky130_fd_sc_hd__o211a_1 _12331_ (.A1(net811),
    .A2(_05191_),
    .B1(_05203_),
    .C1(_05195_),
    .X(_00249_));
 sky130_fd_sc_hd__buf_2 _12332_ (.A(_05177_),
    .X(_05204_));
 sky130_fd_sc_hd__or2_1 _12333_ (.A(net329),
    .B(_05196_),
    .X(_05205_));
 sky130_fd_sc_hd__o211a_1 _12334_ (.A1(net863),
    .A2(_05204_),
    .B1(_05205_),
    .C1(_05195_),
    .X(_00250_));
 sky130_fd_sc_hd__or2_1 _12335_ (.A(net292),
    .B(_05196_),
    .X(_05206_));
 sky130_fd_sc_hd__o211a_1 _12336_ (.A1(net678),
    .A2(_05204_),
    .B1(_05206_),
    .C1(_05195_),
    .X(_00251_));
 sky130_fd_sc_hd__or2_1 _12337_ (.A(net298),
    .B(_05196_),
    .X(_05207_));
 sky130_fd_sc_hd__buf_2 _12338_ (.A(_05127_),
    .X(_05208_));
 sky130_fd_sc_hd__o211a_1 _12339_ (.A1(net540),
    .A2(_05204_),
    .B1(_05207_),
    .C1(_05208_),
    .X(_00252_));
 sky130_fd_sc_hd__clkbuf_2 _12340_ (.A(_05142_),
    .X(_05209_));
 sky130_fd_sc_hd__or2_1 _12341_ (.A(net333),
    .B(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__o211a_1 _12342_ (.A1(net650),
    .A2(_05204_),
    .B1(_05210_),
    .C1(_05208_),
    .X(_00253_));
 sky130_fd_sc_hd__or2_1 _12343_ (.A(net321),
    .B(_05209_),
    .X(_05211_));
 sky130_fd_sc_hd__o211a_1 _12344_ (.A1(net726),
    .A2(_05204_),
    .B1(_05211_),
    .C1(_05208_),
    .X(_00254_));
 sky130_fd_sc_hd__or2_1 _12345_ (.A(net286),
    .B(_05209_),
    .X(_05212_));
 sky130_fd_sc_hd__o211a_1 _12346_ (.A1(net698),
    .A2(_05204_),
    .B1(_05212_),
    .C1(_05208_),
    .X(_00255_));
 sky130_fd_sc_hd__or2_1 _12347_ (.A(net276),
    .B(_05209_),
    .X(_05213_));
 sky130_fd_sc_hd__o211a_1 _12348_ (.A1(net879),
    .A2(_05204_),
    .B1(_05213_),
    .C1(_05208_),
    .X(_00256_));
 sky130_fd_sc_hd__or2_1 _12349_ (.A(net288),
    .B(_05209_),
    .X(_05214_));
 sky130_fd_sc_hd__o211a_1 _12350_ (.A1(net747),
    .A2(_05204_),
    .B1(_05214_),
    .C1(_05208_),
    .X(_00257_));
 sky130_fd_sc_hd__or2_1 _12351_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][27] ),
    .B(_05209_),
    .X(_05215_));
 sky130_fd_sc_hd__o211a_1 _12352_ (.A1(net306),
    .A2(_05204_),
    .B1(_05215_),
    .C1(_05208_),
    .X(_00258_));
 sky130_fd_sc_hd__or2_1 _12353_ (.A(net680),
    .B(_05209_),
    .X(_05216_));
 sky130_fd_sc_hd__o211a_1 _12354_ (.A1(net691),
    .A2(_05204_),
    .B1(_05216_),
    .C1(_05208_),
    .X(_00259_));
 sky130_fd_sc_hd__clkbuf_4 _12355_ (.A(_05177_),
    .X(_05217_));
 sky130_fd_sc_hd__or2_1 _12356_ (.A(net304),
    .B(_05209_),
    .X(_05218_));
 sky130_fd_sc_hd__o211a_1 _12357_ (.A1(net695),
    .A2(_05217_),
    .B1(_05218_),
    .C1(_05208_),
    .X(_00260_));
 sky130_fd_sc_hd__or2_1 _12358_ (.A(net335),
    .B(_05209_),
    .X(_05219_));
 sky130_fd_sc_hd__o211a_1 _12359_ (.A1(net664),
    .A2(_05217_),
    .B1(_05219_),
    .C1(_05208_),
    .X(_00261_));
 sky130_fd_sc_hd__or2_1 _12360_ (.A(net300),
    .B(_05209_),
    .X(_05220_));
 sky130_fd_sc_hd__clkbuf_4 _12361_ (.A(_05127_),
    .X(_05221_));
 sky130_fd_sc_hd__o211a_1 _12362_ (.A1(net929),
    .A2(_05217_),
    .B1(_05220_),
    .C1(_05221_),
    .X(_00262_));
 sky130_fd_sc_hd__clkbuf_2 _12363_ (.A(_05142_),
    .X(_05222_));
 sky130_fd_sc_hd__or2_1 _12364_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][0] ),
    .B(_05222_),
    .X(_05223_));
 sky130_fd_sc_hd__o211a_1 _12365_ (.A1(net495),
    .A2(_05217_),
    .B1(_05223_),
    .C1(_05221_),
    .X(_00263_));
 sky130_fd_sc_hd__or2_1 _12366_ (.A(net432),
    .B(_05222_),
    .X(_05224_));
 sky130_fd_sc_hd__o211a_1 _12367_ (.A1(net466),
    .A2(_05217_),
    .B1(_05224_),
    .C1(_05221_),
    .X(_00264_));
 sky130_fd_sc_hd__or2_1 _12368_ (.A(net835),
    .B(_05222_),
    .X(_05225_));
 sky130_fd_sc_hd__o211a_1 _12369_ (.A1(net848),
    .A2(_05217_),
    .B1(_05225_),
    .C1(_05221_),
    .X(_00265_));
 sky130_fd_sc_hd__or2_1 _12370_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][3] ),
    .B(_05222_),
    .X(_05226_));
 sky130_fd_sc_hd__o211a_1 _12371_ (.A1(net456),
    .A2(_05217_),
    .B1(_05226_),
    .C1(_05221_),
    .X(_00266_));
 sky130_fd_sc_hd__or2_1 _12372_ (.A(net398),
    .B(_05222_),
    .X(_05227_));
 sky130_fd_sc_hd__o211a_1 _12373_ (.A1(net912),
    .A2(_05217_),
    .B1(_05227_),
    .C1(_05221_),
    .X(_00267_));
 sky130_fd_sc_hd__or2_1 _12374_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][5] ),
    .B(_05222_),
    .X(_05228_));
 sky130_fd_sc_hd__o211a_1 _12375_ (.A1(net452),
    .A2(_05217_),
    .B1(_05228_),
    .C1(_05221_),
    .X(_00268_));
 sky130_fd_sc_hd__or2_1 _12376_ (.A(net402),
    .B(_05222_),
    .X(_05229_));
 sky130_fd_sc_hd__o211a_1 _12377_ (.A1(net896),
    .A2(_05217_),
    .B1(_05229_),
    .C1(_05221_),
    .X(_00269_));
 sky130_fd_sc_hd__buf_2 _12378_ (.A(_05177_),
    .X(_05230_));
 sky130_fd_sc_hd__or2_1 _12379_ (.A(net418),
    .B(_05222_),
    .X(_05231_));
 sky130_fd_sc_hd__o211a_1 _12380_ (.A1(net901),
    .A2(_05230_),
    .B1(_05231_),
    .C1(_05221_),
    .X(_00270_));
 sky130_fd_sc_hd__or2_1 _12381_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][8] ),
    .B(_05222_),
    .X(_05232_));
 sky130_fd_sc_hd__o211a_1 _12382_ (.A1(net568),
    .A2(_05230_),
    .B1(_05232_),
    .C1(_05221_),
    .X(_00271_));
 sky130_fd_sc_hd__or2_1 _12383_ (.A(net373),
    .B(_05222_),
    .X(_05233_));
 sky130_fd_sc_hd__buf_2 _12384_ (.A(_05127_),
    .X(_05234_));
 sky130_fd_sc_hd__o211a_1 _12385_ (.A1(net572),
    .A2(_05230_),
    .B1(_05233_),
    .C1(_05234_),
    .X(_00272_));
 sky130_fd_sc_hd__clkbuf_2 _12386_ (.A(_05142_),
    .X(_05235_));
 sky130_fd_sc_hd__or2_1 _12387_ (.A(net357),
    .B(_05235_),
    .X(_05236_));
 sky130_fd_sc_hd__o211a_1 _12388_ (.A1(net807),
    .A2(_05230_),
    .B1(_05236_),
    .C1(_05234_),
    .X(_00273_));
 sky130_fd_sc_hd__or2_1 _12389_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][11] ),
    .B(_05235_),
    .X(_05237_));
 sky130_fd_sc_hd__o211a_1 _12390_ (.A1(net535),
    .A2(_05230_),
    .B1(_05237_),
    .C1(_05234_),
    .X(_00274_));
 sky130_fd_sc_hd__or2_1 _12391_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][12] ),
    .B(_05235_),
    .X(_05238_));
 sky130_fd_sc_hd__o211a_1 _12392_ (.A1(net449),
    .A2(_05230_),
    .B1(_05238_),
    .C1(_05234_),
    .X(_00275_));
 sky130_fd_sc_hd__or2_1 _12393_ (.A(net566),
    .B(_05235_),
    .X(_05239_));
 sky130_fd_sc_hd__o211a_1 _12394_ (.A1(net567),
    .A2(_05230_),
    .B1(_05239_),
    .C1(_05234_),
    .X(_00276_));
 sky130_fd_sc_hd__or2_1 _12395_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][14] ),
    .B(_05235_),
    .X(_05240_));
 sky130_fd_sc_hd__o211a_1 _12396_ (.A1(net515),
    .A2(_05230_),
    .B1(_05240_),
    .C1(_05234_),
    .X(_00277_));
 sky130_fd_sc_hd__or2_1 _12397_ (.A(net323),
    .B(_05235_),
    .X(_05241_));
 sky130_fd_sc_hd__o211a_1 _12398_ (.A1(net505),
    .A2(_05230_),
    .B1(_05241_),
    .C1(_05234_),
    .X(_00278_));
 sky130_fd_sc_hd__or2_1 _12399_ (.A(net346),
    .B(_05235_),
    .X(_05242_));
 sky130_fd_sc_hd__o211a_1 _12400_ (.A1(net480),
    .A2(_05230_),
    .B1(_05242_),
    .C1(_05234_),
    .X(_00279_));
 sky130_fd_sc_hd__buf_2 _12401_ (.A(_05177_),
    .X(_05243_));
 sky130_fd_sc_hd__or2_1 _12402_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][17] ),
    .B(_05235_),
    .X(_05244_));
 sky130_fd_sc_hd__o211a_1 _12403_ (.A1(net319),
    .A2(_05243_),
    .B1(_05244_),
    .C1(_05234_),
    .X(_00280_));
 sky130_fd_sc_hd__or2_1 _12404_ (.A(net341),
    .B(_05235_),
    .X(_05245_));
 sky130_fd_sc_hd__o211a_1 _12405_ (.A1(net345),
    .A2(_05243_),
    .B1(_05245_),
    .C1(_05234_),
    .X(_00281_));
 sky130_fd_sc_hd__or2_1 _12406_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][19] ),
    .B(_05235_),
    .X(_05246_));
 sky130_fd_sc_hd__buf_2 _12407_ (.A(_05127_),
    .X(_05247_));
 sky130_fd_sc_hd__o211a_1 _12408_ (.A1(net329),
    .A2(_05243_),
    .B1(_05246_),
    .C1(_05247_),
    .X(_00282_));
 sky130_fd_sc_hd__clkbuf_2 _12409_ (.A(_05142_),
    .X(_05248_));
 sky130_fd_sc_hd__or2_1 _12410_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][20] ),
    .B(_05248_),
    .X(_05249_));
 sky130_fd_sc_hd__o211a_1 _12411_ (.A1(net292),
    .A2(_05243_),
    .B1(_05249_),
    .C1(_05247_),
    .X(_00283_));
 sky130_fd_sc_hd__or2_1 _12412_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][21] ),
    .B(_05248_),
    .X(_05250_));
 sky130_fd_sc_hd__o211a_1 _12413_ (.A1(net298),
    .A2(_05243_),
    .B1(_05250_),
    .C1(_05247_),
    .X(_00284_));
 sky130_fd_sc_hd__or2_1 _12414_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][22] ),
    .B(_05248_),
    .X(_05251_));
 sky130_fd_sc_hd__o211a_1 _12415_ (.A1(net333),
    .A2(_05243_),
    .B1(_05251_),
    .C1(_05247_),
    .X(_00285_));
 sky130_fd_sc_hd__or2_1 _12416_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][23] ),
    .B(_05248_),
    .X(_05252_));
 sky130_fd_sc_hd__o211a_1 _12417_ (.A1(net321),
    .A2(_05243_),
    .B1(_05252_),
    .C1(_05247_),
    .X(_00286_));
 sky130_fd_sc_hd__or2_1 _12418_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][24] ),
    .B(_05248_),
    .X(_05253_));
 sky130_fd_sc_hd__o211a_1 _12419_ (.A1(net286),
    .A2(_05243_),
    .B1(_05253_),
    .C1(_05247_),
    .X(_00287_));
 sky130_fd_sc_hd__or2_1 _12420_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][25] ),
    .B(_05248_),
    .X(_05254_));
 sky130_fd_sc_hd__o211a_1 _12421_ (.A1(net276),
    .A2(_05243_),
    .B1(_05254_),
    .C1(_05247_),
    .X(_00288_));
 sky130_fd_sc_hd__or2_1 _12422_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][26] ),
    .B(_05248_),
    .X(_05255_));
 sky130_fd_sc_hd__o211a_1 _12423_ (.A1(net288),
    .A2(_05243_),
    .B1(_05255_),
    .C1(_05247_),
    .X(_00289_));
 sky130_fd_sc_hd__clkbuf_8 _12424_ (.A(_05177_),
    .X(_05256_));
 sky130_fd_sc_hd__or2_1 _12425_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][27] ),
    .B(_05248_),
    .X(_05257_));
 sky130_fd_sc_hd__o211a_1 _12426_ (.A1(net369),
    .A2(_05256_),
    .B1(_05257_),
    .C1(_05247_),
    .X(_00290_));
 sky130_fd_sc_hd__or2_1 _12427_ (.A(net308),
    .B(_05248_),
    .X(_05258_));
 sky130_fd_sc_hd__o211a_1 _12428_ (.A1(net680),
    .A2(_05256_),
    .B1(_05258_),
    .C1(_05247_),
    .X(_00291_));
 sky130_fd_sc_hd__or2_1 _12429_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][29] ),
    .B(_05248_),
    .X(_05259_));
 sky130_fd_sc_hd__clkbuf_8 _12430_ (.A(_04868_),
    .X(_05260_));
 sky130_fd_sc_hd__buf_6 _12431_ (.A(_05260_),
    .X(_05261_));
 sky130_fd_sc_hd__o211a_1 _12432_ (.A1(net304),
    .A2(_05256_),
    .B1(_05259_),
    .C1(_05261_),
    .X(_00292_));
 sky130_fd_sc_hd__buf_4 _12433_ (.A(_05142_),
    .X(_05262_));
 sky130_fd_sc_hd__or2_1 _12434_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][30] ),
    .B(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__o211a_1 _12435_ (.A1(net335),
    .A2(_05256_),
    .B1(_05263_),
    .C1(_05261_),
    .X(_00293_));
 sky130_fd_sc_hd__or2_1 _12436_ (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][31] ),
    .B(_05262_),
    .X(_05264_));
 sky130_fd_sc_hd__o211a_1 _12437_ (.A1(net300),
    .A2(_05256_),
    .B1(_05264_),
    .C1(_05261_),
    .X(_00294_));
 sky130_fd_sc_hd__buf_8 _12438_ (.A(net34),
    .X(_05265_));
 sky130_fd_sc_hd__buf_6 _12439_ (.A(net186),
    .X(_05266_));
 sky130_fd_sc_hd__clkbuf_8 _12440_ (.A(net211),
    .X(_05267_));
 sky130_fd_sc_hd__nand2_1 _12441_ (.A(_05267_),
    .B(_04863_),
    .Y(_05268_));
 sky130_fd_sc_hd__buf_6 _12442_ (.A(_05268_),
    .X(_05269_));
 sky130_fd_sc_hd__buf_8 _12443_ (.A(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__mux2_2 _12444_ (.A0(\top_inst.skew_buff_inst.row[0].output_reg[0] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[0] ),
    .S(net211),
    .X(_05271_));
 sky130_fd_sc_hd__clkbuf_4 _12445_ (.A(_05271_),
    .X(_05272_));
 sky130_fd_sc_hd__clkbuf_4 _12446_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[0] ),
    .X(_05273_));
 sky130_fd_sc_hd__and3_1 _12447_ (.A(\top_inst.axis_in_inst.inbuf_valid ),
    .B(_05267_),
    .C(_04857_),
    .X(_05274_));
 sky130_fd_sc_hd__clkbuf_8 _12448_ (.A(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__buf_4 _12449_ (.A(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__or2_1 _12450_ (.A(_05273_),
    .B(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__o211a_1 _12451_ (.A1(_05270_),
    .A2(_05272_),
    .B1(_05277_),
    .C1(_05261_),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_2 _12452_ (.A0(\top_inst.skew_buff_inst.row[0].output_reg[1] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[1] ),
    .S(net211),
    .X(_05278_));
 sky130_fd_sc_hd__clkbuf_4 _12453_ (.A(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__clkbuf_4 _12454_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[1] ),
    .X(_05280_));
 sky130_fd_sc_hd__or2_1 _12455_ (.A(_05280_),
    .B(_05276_),
    .X(_05281_));
 sky130_fd_sc_hd__o211a_1 _12456_ (.A1(_05270_),
    .A2(_05279_),
    .B1(_05281_),
    .C1(_05261_),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_4 _12457_ (.A0(\top_inst.skew_buff_inst.row[0].output_reg[2] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[2] ),
    .S(net213),
    .X(_05282_));
 sky130_fd_sc_hd__buf_2 _12458_ (.A(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__clkbuf_4 _12459_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[2] ),
    .X(_05284_));
 sky130_fd_sc_hd__or2_1 _12460_ (.A(_05284_),
    .B(_05276_),
    .X(_05285_));
 sky130_fd_sc_hd__o211a_1 _12461_ (.A1(_05270_),
    .A2(_05283_),
    .B1(_05285_),
    .C1(_05261_),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_4 _12462_ (.A0(\top_inst.skew_buff_inst.row[0].output_reg[3] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[3] ),
    .S(net211),
    .X(_05286_));
 sky130_fd_sc_hd__buf_2 _12463_ (.A(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__clkbuf_4 _12464_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[3] ),
    .X(_05288_));
 sky130_fd_sc_hd__or2_1 _12465_ (.A(_05288_),
    .B(_05276_),
    .X(_05289_));
 sky130_fd_sc_hd__o211a_1 _12466_ (.A1(_05270_),
    .A2(_05287_),
    .B1(_05289_),
    .C1(_05261_),
    .X(_00298_));
 sky130_fd_sc_hd__clkbuf_4 _12467_ (.A(_05269_),
    .X(_05290_));
 sky130_fd_sc_hd__mux2_2 _12468_ (.A0(\top_inst.skew_buff_inst.row[0].output_reg[4] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[4] ),
    .S(net211),
    .X(_05291_));
 sky130_fd_sc_hd__clkbuf_4 _12469_ (.A(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__clkbuf_4 _12470_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[4] ),
    .X(_05293_));
 sky130_fd_sc_hd__buf_2 _12471_ (.A(_05275_),
    .X(_05294_));
 sky130_fd_sc_hd__or2_1 _12472_ (.A(_05293_),
    .B(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__o211a_1 _12473_ (.A1(_05290_),
    .A2(_05292_),
    .B1(_05295_),
    .C1(_05261_),
    .X(_00299_));
 sky130_fd_sc_hd__mux2_4 _12474_ (.A0(\top_inst.skew_buff_inst.row[0].output_reg[5] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[5] ),
    .S(net213),
    .X(_05296_));
 sky130_fd_sc_hd__buf_4 _12475_ (.A(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__clkbuf_4 _12476_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[5] ),
    .X(_05298_));
 sky130_fd_sc_hd__or2_1 _12477_ (.A(_05298_),
    .B(_05294_),
    .X(_05299_));
 sky130_fd_sc_hd__o211a_1 _12478_ (.A1(_05290_),
    .A2(_05297_),
    .B1(_05299_),
    .C1(_05261_),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _12479_ (.A0(\top_inst.skew_buff_inst.row[0].output_reg[6] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[6] ),
    .S(_05267_),
    .X(_05300_));
 sky130_fd_sc_hd__clkbuf_4 _12480_ (.A(_05300_),
    .X(_05301_));
 sky130_fd_sc_hd__clkbuf_4 _12481_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[6] ),
    .X(_05302_));
 sky130_fd_sc_hd__or2_1 _12482_ (.A(_05302_),
    .B(_05294_),
    .X(_05303_));
 sky130_fd_sc_hd__o211a_1 _12483_ (.A1(_05290_),
    .A2(_05301_),
    .B1(_05303_),
    .C1(_05261_),
    .X(_00301_));
 sky130_fd_sc_hd__buf_2 _12484_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[7] ),
    .X(_05304_));
 sky130_fd_sc_hd__mux2_4 _12485_ (.A0(\top_inst.skew_buff_inst.row[0].output_reg[7] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[7] ),
    .S(_05267_),
    .X(_05305_));
 sky130_fd_sc_hd__clkbuf_4 _12486_ (.A(_05305_),
    .X(_05306_));
 sky130_fd_sc_hd__or2_1 _12487_ (.A(_05269_),
    .B(_05306_),
    .X(_05307_));
 sky130_fd_sc_hd__buf_4 _12488_ (.A(_05260_),
    .X(_05308_));
 sky130_fd_sc_hd__o211a_1 _12489_ (.A1(_05304_),
    .A2(_05276_),
    .B1(_05307_),
    .C1(_05308_),
    .X(_00302_));
 sky130_fd_sc_hd__or2_4 _12490_ (.A(_05267_),
    .B(_04856_),
    .X(_05309_));
 sky130_fd_sc_hd__nor2_2 _12491_ (.A(_04861_),
    .B(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__buf_8 _12492_ (.A(_05310_),
    .X(_05311_));
 sky130_fd_sc_hd__buf_8 _12493_ (.A(_05311_),
    .X(_05312_));
 sky130_fd_sc_hd__buf_12 _12494_ (.A(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__buf_4 _12495_ (.A(_05313_),
    .X(_05314_));
 sky130_fd_sc_hd__buf_6 _12496_ (.A(_05310_),
    .X(_05315_));
 sky130_fd_sc_hd__buf_6 _12497_ (.A(_05315_),
    .X(_05316_));
 sky130_fd_sc_hd__clkbuf_16 _12498_ (.A(_05316_),
    .X(_05317_));
 sky130_fd_sc_hd__nand2_1 _12499_ (.A(_05273_),
    .B(_05272_),
    .Y(_05318_));
 sky130_fd_sc_hd__nand2_1 _12500_ (.A(_05317_),
    .B(_05318_),
    .Y(_05319_));
 sky130_fd_sc_hd__o211a_1 _12501_ (.A1(net950),
    .A2(_05314_),
    .B1(_05319_),
    .C1(_05308_),
    .X(_00303_));
 sky130_fd_sc_hd__a22o_1 _12502_ (.A1(_05280_),
    .A2(_05272_),
    .B1(_05279_),
    .B2(_05273_),
    .X(_05320_));
 sky130_fd_sc_hd__nand2_1 _12503_ (.A(_05280_),
    .B(_05279_),
    .Y(_05321_));
 sky130_fd_sc_hd__or2_1 _12504_ (.A(_05318_),
    .B(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__nor2_2 _12505_ (.A(_05267_),
    .B(_04856_),
    .Y(_05323_));
 sky130_fd_sc_hd__nand2_1 _12506_ (.A(\top_inst.axis_in_inst.inbuf_valid ),
    .B(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__clkbuf_16 _12507_ (.A(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__buf_8 _12508_ (.A(_05325_),
    .X(_05326_));
 sky130_fd_sc_hd__clkbuf_16 _12509_ (.A(_05326_),
    .X(_05327_));
 sky130_fd_sc_hd__buf_8 _12510_ (.A(_05327_),
    .X(_05328_));
 sky130_fd_sc_hd__a21o_1 _12511_ (.A1(_05320_),
    .A2(_05322_),
    .B1(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__o211a_1 _12512_ (.A1(net1026),
    .A2(_05314_),
    .B1(_05329_),
    .C1(_05308_),
    .X(_00304_));
 sky130_fd_sc_hd__nand2_1 _12513_ (.A(_05273_),
    .B(_05283_),
    .Y(_05330_));
 sky130_fd_sc_hd__and3_1 _12514_ (.A(_05280_),
    .B(_05279_),
    .C(_05318_),
    .X(_05331_));
 sky130_fd_sc_hd__xnor2_1 _12515_ (.A(_05330_),
    .B(_05331_),
    .Y(_05332_));
 sky130_fd_sc_hd__a21oi_1 _12516_ (.A1(_05284_),
    .A2(_05272_),
    .B1(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__and3_1 _12517_ (.A(_05284_),
    .B(_05272_),
    .C(_05332_),
    .X(_05334_));
 sky130_fd_sc_hd__buf_8 _12518_ (.A(_05311_),
    .X(_05335_));
 sky130_fd_sc_hd__buf_4 _12519_ (.A(_05335_),
    .X(_05336_));
 sky130_fd_sc_hd__o21ai_1 _12520_ (.A1(_05333_),
    .A2(_05334_),
    .B1(_05336_),
    .Y(_05337_));
 sky130_fd_sc_hd__o211a_1 _12521_ (.A1(net1005),
    .A2(_05314_),
    .B1(_05337_),
    .C1(_05308_),
    .X(_00305_));
 sky130_fd_sc_hd__a22oi_1 _12522_ (.A1(_05288_),
    .A2(_05272_),
    .B1(_05279_),
    .B2(_05284_),
    .Y(_05338_));
 sky130_fd_sc_hd__and4_1 _12523_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[3] ),
    .B(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[2] ),
    .C(_05271_),
    .D(_05278_),
    .X(_05339_));
 sky130_fd_sc_hd__nor2_1 _12524_ (.A(_05338_),
    .B(_05339_),
    .Y(_05340_));
 sky130_fd_sc_hd__nand2_1 _12525_ (.A(_05273_),
    .B(_05287_),
    .Y(_05341_));
 sky130_fd_sc_hd__or2_1 _12526_ (.A(_05321_),
    .B(_05330_),
    .X(_05342_));
 sky130_fd_sc_hd__nand3_1 _12527_ (.A(_05280_),
    .B(_05283_),
    .C(_05342_),
    .Y(_05343_));
 sky130_fd_sc_hd__xor2_1 _12528_ (.A(_05341_),
    .B(_05343_),
    .X(_05344_));
 sky130_fd_sc_hd__nand2_1 _12529_ (.A(_05340_),
    .B(_05344_),
    .Y(_05345_));
 sky130_fd_sc_hd__or2_1 _12530_ (.A(_05340_),
    .B(_05344_),
    .X(_05346_));
 sky130_fd_sc_hd__and2_1 _12531_ (.A(_05345_),
    .B(_05346_),
    .X(_05347_));
 sky130_fd_sc_hd__o21bai_1 _12532_ (.A1(_05283_),
    .A2(_05322_),
    .B1_N(_05334_),
    .Y(_05348_));
 sky130_fd_sc_hd__nor2_1 _12533_ (.A(_05347_),
    .B(_05348_),
    .Y(_05349_));
 sky130_fd_sc_hd__and2_1 _12534_ (.A(_05347_),
    .B(_05348_),
    .X(_05350_));
 sky130_fd_sc_hd__o21ai_1 _12535_ (.A1(_05349_),
    .A2(_05350_),
    .B1(_05336_),
    .Y(_05351_));
 sky130_fd_sc_hd__o211a_1 _12536_ (.A1(net1048),
    .A2(_05314_),
    .B1(_05351_),
    .C1(_05308_),
    .X(_00306_));
 sky130_fd_sc_hd__buf_8 _12537_ (.A(_04869_),
    .X(_05352_));
 sky130_fd_sc_hd__buf_6 _12538_ (.A(_05325_),
    .X(_05353_));
 sky130_fd_sc_hd__buf_8 _12539_ (.A(_05353_),
    .X(_05354_));
 sky130_fd_sc_hd__and4_1 _12540_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[1] ),
    .B(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[0] ),
    .C(_05282_),
    .D(_05287_),
    .X(_05355_));
 sky130_fd_sc_hd__nor2_1 _12541_ (.A(_05342_),
    .B(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__inv_2 _12542_ (.A(_05355_),
    .Y(_05357_));
 sky130_fd_sc_hd__and4_1 _12543_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[1] ),
    .B(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[0] ),
    .C(_05286_),
    .D(_05291_),
    .X(_05358_));
 sky130_fd_sc_hd__a22oi_1 _12544_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[1] ),
    .A2(_05286_),
    .B1(_05291_),
    .B2(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[0] ),
    .Y(_05359_));
 sky130_fd_sc_hd__nor2_1 _12545_ (.A(_05358_),
    .B(_05359_),
    .Y(_05360_));
 sky130_fd_sc_hd__xnor2_1 _12546_ (.A(_05339_),
    .B(_05360_),
    .Y(_05361_));
 sky130_fd_sc_hd__xnor2_1 _12547_ (.A(_05357_),
    .B(_05361_),
    .Y(_05362_));
 sky130_fd_sc_hd__and4_1 _12548_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[3] ),
    .C(_05271_),
    .D(_05278_),
    .X(_05363_));
 sky130_fd_sc_hd__a22o_1 _12549_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[4] ),
    .A2(_05271_),
    .B1(_05278_),
    .B2(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[3] ),
    .X(_05364_));
 sky130_fd_sc_hd__and4b_1 _12550_ (.A_N(_05363_),
    .B(_05284_),
    .C(_05283_),
    .D(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__inv_2 _12551_ (.A(_05364_),
    .Y(_05366_));
 sky130_fd_sc_hd__o2bb2a_1 _12552_ (.A1_N(_05284_),
    .A2_N(_05283_),
    .B1(_05363_),
    .B2(_05366_),
    .X(_05367_));
 sky130_fd_sc_hd__nor2_1 _12553_ (.A(_05365_),
    .B(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__xnor2_1 _12554_ (.A(_05362_),
    .B(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__xor2_1 _12555_ (.A(_05345_),
    .B(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__xnor2_1 _12556_ (.A(_05356_),
    .B(_05370_),
    .Y(_05371_));
 sky130_fd_sc_hd__nand2_1 _12557_ (.A(_05350_),
    .B(_05371_),
    .Y(_05372_));
 sky130_fd_sc_hd__o21a_1 _12558_ (.A1(_05350_),
    .A2(_05371_),
    .B1(_05315_),
    .X(_05373_));
 sky130_fd_sc_hd__a22o_1 _12559_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[4] ),
    .A2(_05354_),
    .B1(_05372_),
    .B2(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__and2_1 _12560_ (.A(_05352_),
    .B(_05374_),
    .X(_05375_));
 sky130_fd_sc_hd__clkbuf_1 _12561_ (.A(_05375_),
    .X(_00307_));
 sky130_fd_sc_hd__or3_1 _12562_ (.A(_05362_),
    .B(_05365_),
    .C(_05367_),
    .X(_05376_));
 sky130_fd_sc_hd__nand2_1 _12563_ (.A(_05298_),
    .B(_05272_),
    .Y(_05377_));
 sky130_fd_sc_hd__a22o_1 _12564_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[4] ),
    .A2(_05278_),
    .B1(_05282_),
    .B2(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[3] ),
    .X(_05378_));
 sky130_fd_sc_hd__nand4_1 _12565_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[3] ),
    .C(_05279_),
    .D(_05282_),
    .Y(_05379_));
 sky130_fd_sc_hd__nand2_1 _12566_ (.A(_05378_),
    .B(_05379_),
    .Y(_05380_));
 sky130_fd_sc_hd__and2_1 _12567_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[2] ),
    .B(_05286_),
    .X(_05381_));
 sky130_fd_sc_hd__xor2_1 _12568_ (.A(_05380_),
    .B(_05381_),
    .X(_05382_));
 sky130_fd_sc_hd__xor2_1 _12569_ (.A(_05377_),
    .B(_05382_),
    .X(_05383_));
 sky130_fd_sc_hd__a31o_1 _12570_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[2] ),
    .A2(_05283_),
    .A3(_05364_),
    .B1(_05363_),
    .X(_05384_));
 sky130_fd_sc_hd__and4_1 _12571_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[1] ),
    .B(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[0] ),
    .C(_05291_),
    .D(_05296_),
    .X(_05385_));
 sky130_fd_sc_hd__a22oi_1 _12572_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[1] ),
    .A2(_05292_),
    .B1(_05296_),
    .B2(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[0] ),
    .Y(_05386_));
 sky130_fd_sc_hd__nor2_1 _12573_ (.A(_05385_),
    .B(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__xor2_1 _12574_ (.A(_05384_),
    .B(_05387_),
    .X(_05388_));
 sky130_fd_sc_hd__xnor2_1 _12575_ (.A(_05358_),
    .B(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__xor2_1 _12576_ (.A(_05383_),
    .B(_05389_),
    .X(_05390_));
 sky130_fd_sc_hd__xor2_1 _12577_ (.A(_05376_),
    .B(_05390_),
    .X(_05391_));
 sky130_fd_sc_hd__nor2_1 _12578_ (.A(_05357_),
    .B(_05361_),
    .Y(_05392_));
 sky130_fd_sc_hd__a21o_1 _12579_ (.A1(_05339_),
    .A2(_05360_),
    .B1(_05392_),
    .X(_05393_));
 sky130_fd_sc_hd__xnor2_1 _12580_ (.A(_05391_),
    .B(_05393_),
    .Y(_05394_));
 sky130_fd_sc_hd__or2b_1 _12581_ (.A(_05345_),
    .B_N(_05369_),
    .X(_05395_));
 sky130_fd_sc_hd__o31a_1 _12582_ (.A1(_05342_),
    .A2(_05355_),
    .A3(_05370_),
    .B1(_05395_),
    .X(_05396_));
 sky130_fd_sc_hd__xnor2_1 _12583_ (.A(_05394_),
    .B(_05396_),
    .Y(_05397_));
 sky130_fd_sc_hd__or2_1 _12584_ (.A(_05372_),
    .B(_05397_),
    .X(_05398_));
 sky130_fd_sc_hd__buf_8 _12585_ (.A(_05325_),
    .X(_05399_));
 sky130_fd_sc_hd__a21oi_1 _12586_ (.A1(_05372_),
    .A2(_05397_),
    .B1(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__a22o_1 _12587_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[5] ),
    .A2(_05354_),
    .B1(_05398_),
    .B2(_05400_),
    .X(_05401_));
 sky130_fd_sc_hd__and2_1 _12588_ (.A(_05352_),
    .B(_05401_),
    .X(_05402_));
 sky130_fd_sc_hd__clkbuf_1 _12589_ (.A(_05402_),
    .X(_00308_));
 sky130_fd_sc_hd__buf_8 _12590_ (.A(_05327_),
    .X(_05403_));
 sky130_fd_sc_hd__nand2_1 _12591_ (.A(net982),
    .B(_05403_),
    .Y(_05404_));
 sky130_fd_sc_hd__clkbuf_16 _12592_ (.A(_05325_),
    .X(_05405_));
 sky130_fd_sc_hd__buf_8 _12593_ (.A(_05405_),
    .X(_05406_));
 sky130_fd_sc_hd__or2_1 _12594_ (.A(_05394_),
    .B(_05396_),
    .X(_05407_));
 sky130_fd_sc_hd__or2_1 _12595_ (.A(_05376_),
    .B(_05390_),
    .X(_05408_));
 sky130_fd_sc_hd__nand2_1 _12596_ (.A(_05391_),
    .B(_05393_),
    .Y(_05409_));
 sky130_fd_sc_hd__inv_2 _12597_ (.A(_05389_),
    .Y(_05410_));
 sky130_fd_sc_hd__nand2_1 _12598_ (.A(_05383_),
    .B(_05410_),
    .Y(_05411_));
 sky130_fd_sc_hd__or2_1 _12599_ (.A(_05377_),
    .B(_05382_),
    .X(_05412_));
 sky130_fd_sc_hd__a22o_1 _12600_ (.A1(_05302_),
    .A2(_05272_),
    .B1(_05279_),
    .B2(_05298_),
    .X(_05413_));
 sky130_fd_sc_hd__nand4_2 _12601_ (.A(_05302_),
    .B(_05298_),
    .C(_05272_),
    .D(_05279_),
    .Y(_05414_));
 sky130_fd_sc_hd__nand2_1 _12602_ (.A(_05413_),
    .B(_05414_),
    .Y(_05415_));
 sky130_fd_sc_hd__a22oi_1 _12603_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[4] ),
    .A2(_05282_),
    .B1(_05287_),
    .B2(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[3] ),
    .Y(_05416_));
 sky130_fd_sc_hd__and4_1 _12604_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[3] ),
    .C(_05282_),
    .D(_05287_),
    .X(_05417_));
 sky130_fd_sc_hd__nor2_1 _12605_ (.A(_05416_),
    .B(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__nand2_1 _12606_ (.A(_05284_),
    .B(_05292_),
    .Y(_05419_));
 sky130_fd_sc_hd__xnor2_1 _12607_ (.A(_05418_),
    .B(_05419_),
    .Y(_05420_));
 sky130_fd_sc_hd__xor2_1 _12608_ (.A(_05415_),
    .B(_05420_),
    .X(_05421_));
 sky130_fd_sc_hd__xnor2_1 _12609_ (.A(_05412_),
    .B(_05421_),
    .Y(_05422_));
 sky130_fd_sc_hd__a21bo_1 _12610_ (.A1(_05378_),
    .A2(_05381_),
    .B1_N(_05379_),
    .X(_05423_));
 sky130_fd_sc_hd__and4_1 _12611_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[1] ),
    .B(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[0] ),
    .C(_05296_),
    .D(_05300_),
    .X(_05424_));
 sky130_fd_sc_hd__a22oi_1 _12612_ (.A1(_05280_),
    .A2(_05297_),
    .B1(_05301_),
    .B2(_05273_),
    .Y(_05425_));
 sky130_fd_sc_hd__nor2_1 _12613_ (.A(_05424_),
    .B(_05425_),
    .Y(_05426_));
 sky130_fd_sc_hd__xor2_1 _12614_ (.A(_05423_),
    .B(_05426_),
    .X(_05427_));
 sky130_fd_sc_hd__nor2_1 _12615_ (.A(_05385_),
    .B(_05427_),
    .Y(_05428_));
 sky130_fd_sc_hd__and2_1 _12616_ (.A(_05385_),
    .B(_05427_),
    .X(_05429_));
 sky130_fd_sc_hd__or2_1 _12617_ (.A(_05428_),
    .B(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__xnor2_1 _12618_ (.A(_05422_),
    .B(_05430_),
    .Y(_05431_));
 sky130_fd_sc_hd__xnor2_1 _12619_ (.A(_05411_),
    .B(_05431_),
    .Y(_05432_));
 sky130_fd_sc_hd__a22o_1 _12620_ (.A1(_05384_),
    .A2(_05387_),
    .B1(_05388_),
    .B2(_05358_),
    .X(_05433_));
 sky130_fd_sc_hd__xor2_1 _12621_ (.A(_05432_),
    .B(_05433_),
    .X(_05434_));
 sky130_fd_sc_hd__a21oi_2 _12622_ (.A1(_05408_),
    .A2(_05409_),
    .B1(_05434_),
    .Y(_05435_));
 sky130_fd_sc_hd__and3_1 _12623_ (.A(_05408_),
    .B(_05409_),
    .C(_05434_),
    .X(_05436_));
 sky130_fd_sc_hd__a211oi_2 _12624_ (.A1(_05407_),
    .A2(_05398_),
    .B1(_05435_),
    .C1(_05436_),
    .Y(_05437_));
 sky130_fd_sc_hd__o211a_1 _12625_ (.A1(_05435_),
    .A2(_05436_),
    .B1(_05407_),
    .C1(_05398_),
    .X(_05438_));
 sky130_fd_sc_hd__or3_1 _12626_ (.A(_05406_),
    .B(_05437_),
    .C(_05438_),
    .X(_05439_));
 sky130_fd_sc_hd__buf_8 _12627_ (.A(_04867_),
    .X(_05440_));
 sky130_fd_sc_hd__a21oi_1 _12628_ (.A1(_05404_),
    .A2(_05439_),
    .B1(_05440_),
    .Y(_00309_));
 sky130_fd_sc_hd__nor2_1 _12629_ (.A(_05411_),
    .B(_05431_),
    .Y(_05441_));
 sky130_fd_sc_hd__and2b_1 _12630_ (.A_N(_05432_),
    .B(_05433_),
    .X(_05442_));
 sky130_fd_sc_hd__and2_1 _12631_ (.A(_05423_),
    .B(_05426_),
    .X(_05443_));
 sky130_fd_sc_hd__or2_1 _12632_ (.A(_05412_),
    .B(_05421_),
    .X(_05444_));
 sky130_fd_sc_hd__or2_1 _12633_ (.A(_05422_),
    .B(_05430_),
    .X(_05445_));
 sky130_fd_sc_hd__and3_1 _12634_ (.A(_05413_),
    .B(_05414_),
    .C(_05420_),
    .X(_05446_));
 sky130_fd_sc_hd__inv_2 _12635_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[7] ),
    .Y(_05447_));
 sky130_fd_sc_hd__a2bb2o_1 _12636_ (.A1_N(_05447_),
    .A2_N(_05271_),
    .B1(_05279_),
    .B2(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[6] ),
    .X(_05448_));
 sky130_fd_sc_hd__inv_2 _12637_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[6] ),
    .Y(_05449_));
 sky130_fd_sc_hd__or4b_1 _12638_ (.A(_05447_),
    .B(_05449_),
    .C(_05271_),
    .D_N(_05278_),
    .X(_05450_));
 sky130_fd_sc_hd__nand2_1 _12639_ (.A(_05448_),
    .B(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__and2_1 _12640_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[5] ),
    .B(_05283_),
    .X(_05452_));
 sky130_fd_sc_hd__xor2_1 _12641_ (.A(_05451_),
    .B(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__xnor2_1 _12642_ (.A(_05414_),
    .B(_05453_),
    .Y(_05454_));
 sky130_fd_sc_hd__a22oi_1 _12643_ (.A1(_05293_),
    .A2(_05287_),
    .B1(_05292_),
    .B2(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[3] ),
    .Y(_05455_));
 sky130_fd_sc_hd__and4_1 _12644_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[3] ),
    .C(_05287_),
    .D(_05291_),
    .X(_05456_));
 sky130_fd_sc_hd__or2_1 _12645_ (.A(_05455_),
    .B(_05456_),
    .X(_05457_));
 sky130_fd_sc_hd__nand2_1 _12646_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[2] ),
    .B(_05297_),
    .Y(_05458_));
 sky130_fd_sc_hd__xnor2_1 _12647_ (.A(_05457_),
    .B(_05458_),
    .Y(_05459_));
 sky130_fd_sc_hd__xor2_1 _12648_ (.A(_05454_),
    .B(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__xnor2_1 _12649_ (.A(_05446_),
    .B(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__a31o_1 _12650_ (.A1(_05284_),
    .A2(_05292_),
    .A3(_05418_),
    .B1(_05417_),
    .X(_05462_));
 sky130_fd_sc_hd__a22o_1 _12651_ (.A1(_05280_),
    .A2(_05301_),
    .B1(_05305_),
    .B2(_05273_),
    .X(_05463_));
 sky130_fd_sc_hd__and4_1 _12652_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[1] ),
    .B(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[0] ),
    .C(_05300_),
    .D(_05305_),
    .X(_05464_));
 sky130_fd_sc_hd__inv_2 _12653_ (.A(_05464_),
    .Y(_05465_));
 sky130_fd_sc_hd__and3_1 _12654_ (.A(_05304_),
    .B(_05463_),
    .C(_05465_),
    .X(_05466_));
 sky130_fd_sc_hd__a21oi_1 _12655_ (.A1(_05463_),
    .A2(_05465_),
    .B1(_05304_),
    .Y(_05467_));
 sky130_fd_sc_hd__or2_1 _12656_ (.A(_05466_),
    .B(_05467_),
    .X(_05468_));
 sky130_fd_sc_hd__xnor2_1 _12657_ (.A(_05462_),
    .B(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__xnor2_1 _12658_ (.A(_05424_),
    .B(_05469_),
    .Y(_05470_));
 sky130_fd_sc_hd__xnor2_1 _12659_ (.A(_05461_),
    .B(_05470_),
    .Y(_05471_));
 sky130_fd_sc_hd__a21o_2 _12660_ (.A1(_05444_),
    .A2(_05445_),
    .B1(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__nand3_2 _12661_ (.A(_05444_),
    .B(_05445_),
    .C(_05471_),
    .Y(_05473_));
 sky130_fd_sc_hd__o211ai_4 _12662_ (.A1(_05443_),
    .A2(_05429_),
    .B1(_05472_),
    .C1(_05473_),
    .Y(_05474_));
 sky130_fd_sc_hd__a211o_1 _12663_ (.A1(_05472_),
    .A2(_05473_),
    .B1(_05443_),
    .C1(_05429_),
    .X(_05475_));
 sky130_fd_sc_hd__o211ai_4 _12664_ (.A1(_05441_),
    .A2(_05442_),
    .B1(_05474_),
    .C1(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__a211o_1 _12665_ (.A1(_05474_),
    .A2(_05475_),
    .B1(_05441_),
    .C1(_05442_),
    .X(_05477_));
 sky130_fd_sc_hd__a211o_1 _12666_ (.A1(_05476_),
    .A2(_05477_),
    .B1(_05435_),
    .C1(_05437_),
    .X(_05478_));
 sky130_fd_sc_hd__o211ai_2 _12667_ (.A1(_05435_),
    .A2(_05437_),
    .B1(_05476_),
    .C1(_05477_),
    .Y(_05479_));
 sky130_fd_sc_hd__and2_1 _12668_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[7] ),
    .B(_05326_),
    .X(_05480_));
 sky130_fd_sc_hd__a31o_1 _12669_ (.A1(_05335_),
    .A2(_05478_),
    .A3(_05479_),
    .B1(_05480_),
    .X(_05481_));
 sky130_fd_sc_hd__and2_1 _12670_ (.A(_05352_),
    .B(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__clkbuf_1 _12671_ (.A(_05482_),
    .X(_00310_));
 sky130_fd_sc_hd__nand2_1 _12672_ (.A(net1013),
    .B(_05403_),
    .Y(_05483_));
 sky130_fd_sc_hd__or2b_1 _12673_ (.A(_05468_),
    .B_N(_05462_),
    .X(_05484_));
 sky130_fd_sc_hd__nand2_1 _12674_ (.A(_05424_),
    .B(_05469_),
    .Y(_05485_));
 sky130_fd_sc_hd__nand2_1 _12675_ (.A(_05446_),
    .B(_05460_),
    .Y(_05486_));
 sky130_fd_sc_hd__or2_1 _12676_ (.A(_05461_),
    .B(_05470_),
    .X(_05487_));
 sky130_fd_sc_hd__inv_2 _12677_ (.A(_05278_),
    .Y(_05488_));
 sky130_fd_sc_hd__a22o_1 _12678_ (.A1(_05304_),
    .A2(_05488_),
    .B1(_05283_),
    .B2(_05302_),
    .X(_05489_));
 sky130_fd_sc_hd__inv_2 _12679_ (.A(_05282_),
    .Y(_05490_));
 sky130_fd_sc_hd__or4_1 _12680_ (.A(_05447_),
    .B(_05449_),
    .C(_05279_),
    .D(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__nand2_1 _12681_ (.A(_05489_),
    .B(_05491_),
    .Y(_05492_));
 sky130_fd_sc_hd__nand2_1 _12682_ (.A(_05298_),
    .B(_05287_),
    .Y(_05493_));
 sky130_fd_sc_hd__xnor2_2 _12683_ (.A(_05492_),
    .B(_05493_),
    .Y(_05494_));
 sky130_fd_sc_hd__a21boi_2 _12684_ (.A1(_05448_),
    .A2(_05452_),
    .B1_N(_05450_),
    .Y(_05495_));
 sky130_fd_sc_hd__xnor2_2 _12685_ (.A(_05494_),
    .B(_05495_),
    .Y(_05496_));
 sky130_fd_sc_hd__a22oi_2 _12686_ (.A1(_05293_),
    .A2(_05292_),
    .B1(_05297_),
    .B2(_05288_),
    .Y(_05497_));
 sky130_fd_sc_hd__and4_1 _12687_ (.A(_05293_),
    .B(_05288_),
    .C(_05292_),
    .D(_05297_),
    .X(_05498_));
 sky130_fd_sc_hd__or2_1 _12688_ (.A(_05497_),
    .B(_05498_),
    .X(_05499_));
 sky130_fd_sc_hd__nand2_1 _12689_ (.A(_05284_),
    .B(_05301_),
    .Y(_05500_));
 sky130_fd_sc_hd__xnor2_2 _12690_ (.A(_05499_),
    .B(_05500_),
    .Y(_05501_));
 sky130_fd_sc_hd__xnor2_2 _12691_ (.A(_05496_),
    .B(_05501_),
    .Y(_05502_));
 sky130_fd_sc_hd__or2_1 _12692_ (.A(_05414_),
    .B(_05453_),
    .X(_05503_));
 sky130_fd_sc_hd__o21a_1 _12693_ (.A1(_05454_),
    .A2(_05459_),
    .B1(_05503_),
    .X(_05504_));
 sky130_fd_sc_hd__xor2_2 _12694_ (.A(_05502_),
    .B(_05504_),
    .X(_05505_));
 sky130_fd_sc_hd__o21ba_1 _12695_ (.A1(_05455_),
    .A2(_05458_),
    .B1_N(_05456_),
    .X(_05506_));
 sky130_fd_sc_hd__o21ai_4 _12696_ (.A1(_05280_),
    .A2(_05273_),
    .B1(_05305_),
    .Y(_05507_));
 sky130_fd_sc_hd__and3_1 _12697_ (.A(_05280_),
    .B(_05273_),
    .C(_05305_),
    .X(_05508_));
 sky130_fd_sc_hd__or3_4 _12698_ (.A(_05506_),
    .B(_05507_),
    .C(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__o21ai_1 _12699_ (.A1(_05507_),
    .A2(_05508_),
    .B1(_05506_),
    .Y(_05510_));
 sky130_fd_sc_hd__and2_1 _12700_ (.A(_05509_),
    .B(_05510_),
    .X(_05511_));
 sky130_fd_sc_hd__o21ai_2 _12701_ (.A1(_05464_),
    .A2(_05466_),
    .B1(_05511_),
    .Y(_05512_));
 sky130_fd_sc_hd__or3_1 _12702_ (.A(_05464_),
    .B(_05466_),
    .C(_05511_),
    .X(_05513_));
 sky130_fd_sc_hd__and2_1 _12703_ (.A(_05512_),
    .B(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__xnor2_2 _12704_ (.A(_05505_),
    .B(_05514_),
    .Y(_05515_));
 sky130_fd_sc_hd__a21oi_4 _12705_ (.A1(_05486_),
    .A2(_05487_),
    .B1(_05515_),
    .Y(_05516_));
 sky130_fd_sc_hd__and3_1 _12706_ (.A(_05486_),
    .B(_05487_),
    .C(_05515_),
    .X(_05517_));
 sky130_fd_sc_hd__a211oi_4 _12707_ (.A1(_05484_),
    .A2(_05485_),
    .B1(_05516_),
    .C1(_05517_),
    .Y(_05518_));
 sky130_fd_sc_hd__o211a_1 _12708_ (.A1(_05516_),
    .A2(_05517_),
    .B1(_05484_),
    .C1(_05485_),
    .X(_05519_));
 sky130_fd_sc_hd__a211oi_4 _12709_ (.A1(_05472_),
    .A2(_05474_),
    .B1(_05518_),
    .C1(_05519_),
    .Y(_05520_));
 sky130_fd_sc_hd__o211a_1 _12710_ (.A1(_05518_),
    .A2(_05519_),
    .B1(_05472_),
    .C1(_05474_),
    .X(_05521_));
 sky130_fd_sc_hd__a211oi_2 _12711_ (.A1(_05476_),
    .A2(_05479_),
    .B1(_05520_),
    .C1(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__o211a_1 _12712_ (.A1(_05520_),
    .A2(_05521_),
    .B1(_05476_),
    .C1(_05479_),
    .X(_05523_));
 sky130_fd_sc_hd__or3_1 _12713_ (.A(_05406_),
    .B(_05522_),
    .C(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__a21oi_1 _12714_ (.A1(_05483_),
    .A2(_05524_),
    .B1(_05440_),
    .Y(_00311_));
 sky130_fd_sc_hd__or2_1 _12715_ (.A(_05502_),
    .B(_05504_),
    .X(_05525_));
 sky130_fd_sc_hd__nand2_1 _12716_ (.A(_05505_),
    .B(_05514_),
    .Y(_05526_));
 sky130_fd_sc_hd__a22o_1 _12717_ (.A1(_05304_),
    .A2(_05490_),
    .B1(_05287_),
    .B2(_05302_),
    .X(_05527_));
 sky130_fd_sc_hd__inv_2 _12718_ (.A(_05286_),
    .Y(_05528_));
 sky130_fd_sc_hd__or4_1 _12719_ (.A(_05447_),
    .B(_05449_),
    .C(_05283_),
    .D(_05528_),
    .X(_05529_));
 sky130_fd_sc_hd__nand2_1 _12720_ (.A(_05527_),
    .B(_05529_),
    .Y(_05530_));
 sky130_fd_sc_hd__nand2_1 _12721_ (.A(_05298_),
    .B(_05292_),
    .Y(_05531_));
 sky130_fd_sc_hd__xnor2_1 _12722_ (.A(_05530_),
    .B(_05531_),
    .Y(_05532_));
 sky130_fd_sc_hd__o21a_1 _12723_ (.A1(_05492_),
    .A2(_05493_),
    .B1(_05491_),
    .X(_05533_));
 sky130_fd_sc_hd__xnor2_1 _12724_ (.A(_05532_),
    .B(_05533_),
    .Y(_05534_));
 sky130_fd_sc_hd__a22oi_2 _12725_ (.A1(_05293_),
    .A2(_05297_),
    .B1(_05301_),
    .B2(_05288_),
    .Y(_05535_));
 sky130_fd_sc_hd__and4_1 _12726_ (.A(_05293_),
    .B(_05288_),
    .C(_05297_),
    .D(_05301_),
    .X(_05536_));
 sky130_fd_sc_hd__nor2_1 _12727_ (.A(_05535_),
    .B(_05536_),
    .Y(_05537_));
 sky130_fd_sc_hd__nand2_2 _12728_ (.A(_05284_),
    .B(_05306_),
    .Y(_05538_));
 sky130_fd_sc_hd__xor2_1 _12729_ (.A(_05537_),
    .B(_05538_),
    .X(_05539_));
 sky130_fd_sc_hd__or2_1 _12730_ (.A(_05534_),
    .B(_05539_),
    .X(_05540_));
 sky130_fd_sc_hd__nand2_1 _12731_ (.A(_05534_),
    .B(_05539_),
    .Y(_05541_));
 sky130_fd_sc_hd__nand2_1 _12732_ (.A(_05540_),
    .B(_05541_),
    .Y(_05542_));
 sky130_fd_sc_hd__or2_1 _12733_ (.A(_05494_),
    .B(_05495_),
    .X(_05543_));
 sky130_fd_sc_hd__o21a_1 _12734_ (.A1(_05496_),
    .A2(_05501_),
    .B1(_05543_),
    .X(_05544_));
 sky130_fd_sc_hd__xor2_1 _12735_ (.A(_05542_),
    .B(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__o21ba_1 _12736_ (.A1(_05497_),
    .A2(_05500_),
    .B1_N(_05498_),
    .X(_05546_));
 sky130_fd_sc_hd__or2_1 _12737_ (.A(_05507_),
    .B(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__nand2_1 _12738_ (.A(_05507_),
    .B(_05546_),
    .Y(_05548_));
 sky130_fd_sc_hd__and2_1 _12739_ (.A(_05547_),
    .B(_05548_),
    .X(_05549_));
 sky130_fd_sc_hd__and2_2 _12740_ (.A(_05545_),
    .B(_05549_),
    .X(_05550_));
 sky130_fd_sc_hd__nor2_1 _12741_ (.A(_05545_),
    .B(_05549_),
    .Y(_05551_));
 sky130_fd_sc_hd__a211oi_4 _12742_ (.A1(_05525_),
    .A2(_05526_),
    .B1(_05550_),
    .C1(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__o211a_1 _12743_ (.A1(_05550_),
    .A2(_05551_),
    .B1(_05525_),
    .C1(_05526_),
    .X(_05553_));
 sky130_fd_sc_hd__a211o_2 _12744_ (.A1(_05509_),
    .A2(_05512_),
    .B1(_05552_),
    .C1(_05553_),
    .X(_05554_));
 sky130_fd_sc_hd__o211ai_4 _12745_ (.A1(_05552_),
    .A2(_05553_),
    .B1(_05509_),
    .C1(_05512_),
    .Y(_05555_));
 sky130_fd_sc_hd__o211ai_4 _12746_ (.A1(_05516_),
    .A2(_05518_),
    .B1(_05554_),
    .C1(_05555_),
    .Y(_05556_));
 sky130_fd_sc_hd__a211o_1 _12747_ (.A1(_05554_),
    .A2(_05555_),
    .B1(_05516_),
    .C1(_05518_),
    .X(_05557_));
 sky130_fd_sc_hd__o211ai_2 _12748_ (.A1(_05520_),
    .A2(_05522_),
    .B1(_05556_),
    .C1(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__a211o_1 _12749_ (.A1(_05556_),
    .A2(_05557_),
    .B1(_05520_),
    .C1(_05522_),
    .X(_05559_));
 sky130_fd_sc_hd__a21o_1 _12750_ (.A1(_05558_),
    .A2(_05559_),
    .B1(_05328_),
    .X(_05560_));
 sky130_fd_sc_hd__o211a_1 _12751_ (.A1(net1084),
    .A2(_05314_),
    .B1(_05560_),
    .C1(_05308_),
    .X(_00312_));
 sky130_fd_sc_hd__nand2_1 _12752_ (.A(net1010),
    .B(_05403_),
    .Y(_05561_));
 sky130_fd_sc_hd__inv_2 _12753_ (.A(_05552_),
    .Y(_05562_));
 sky130_fd_sc_hd__nor2_1 _12754_ (.A(_05542_),
    .B(_05544_),
    .Y(_05563_));
 sky130_fd_sc_hd__or2_1 _12755_ (.A(_05532_),
    .B(_05533_),
    .X(_05564_));
 sky130_fd_sc_hd__a22o_1 _12756_ (.A1(_05304_),
    .A2(_05528_),
    .B1(_05292_),
    .B2(_05302_),
    .X(_05565_));
 sky130_fd_sc_hd__and2b_1 _12757_ (.A_N(_05267_),
    .B(\top_inst.skew_buff_inst.row[0].output_reg[4] ),
    .X(_05566_));
 sky130_fd_sc_hd__a21oi_2 _12758_ (.A1(\top_inst.axis_in_inst.inbuf_bus[4] ),
    .A2(_05267_),
    .B1(_05566_),
    .Y(_05567_));
 sky130_fd_sc_hd__or4_1 _12759_ (.A(_05447_),
    .B(_05449_),
    .C(_05287_),
    .D(_05567_),
    .X(_05568_));
 sky130_fd_sc_hd__nand2_1 _12760_ (.A(_05565_),
    .B(_05568_),
    .Y(_05569_));
 sky130_fd_sc_hd__nand2_1 _12761_ (.A(_05298_),
    .B(_05297_),
    .Y(_05570_));
 sky130_fd_sc_hd__xnor2_2 _12762_ (.A(_05569_),
    .B(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__o21a_1 _12763_ (.A1(_05530_),
    .A2(_05531_),
    .B1(_05529_),
    .X(_05572_));
 sky130_fd_sc_hd__xnor2_1 _12764_ (.A(_05571_),
    .B(_05572_),
    .Y(_05573_));
 sky130_fd_sc_hd__a22oi_2 _12765_ (.A1(_05293_),
    .A2(_05301_),
    .B1(_05306_),
    .B2(_05288_),
    .Y(_05574_));
 sky130_fd_sc_hd__and4_1 _12766_ (.A(_05293_),
    .B(_05288_),
    .C(_05301_),
    .D(_05306_),
    .X(_05575_));
 sky130_fd_sc_hd__nor2_1 _12767_ (.A(_05574_),
    .B(_05575_),
    .Y(_05576_));
 sky130_fd_sc_hd__xnor2_1 _12768_ (.A(_05538_),
    .B(_05576_),
    .Y(_05577_));
 sky130_fd_sc_hd__xor2_1 _12769_ (.A(_05573_),
    .B(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__a21o_1 _12770_ (.A1(_05564_),
    .A2(_05540_),
    .B1(_05578_),
    .X(_05579_));
 sky130_fd_sc_hd__nand3_1 _12771_ (.A(_05564_),
    .B(_05540_),
    .C(_05578_),
    .Y(_05580_));
 sky130_fd_sc_hd__o21ba_1 _12772_ (.A1(_05535_),
    .A2(_05538_),
    .B1_N(_05536_),
    .X(_05581_));
 sky130_fd_sc_hd__or2_1 _12773_ (.A(_05507_),
    .B(_05581_),
    .X(_05582_));
 sky130_fd_sc_hd__nand2_1 _12774_ (.A(_05507_),
    .B(_05581_),
    .Y(_05583_));
 sky130_fd_sc_hd__and2_1 _12775_ (.A(_05582_),
    .B(_05583_),
    .X(_05584_));
 sky130_fd_sc_hd__nand3_1 _12776_ (.A(_05579_),
    .B(_05580_),
    .C(_05584_),
    .Y(_05585_));
 sky130_fd_sc_hd__a21o_1 _12777_ (.A1(_05579_),
    .A2(_05580_),
    .B1(_05584_),
    .X(_05586_));
 sky130_fd_sc_hd__o211ai_1 _12778_ (.A1(_05563_),
    .A2(_05550_),
    .B1(_05585_),
    .C1(_05586_),
    .Y(_05587_));
 sky130_fd_sc_hd__a211o_1 _12779_ (.A1(_05585_),
    .A2(_05586_),
    .B1(_05563_),
    .C1(_05550_),
    .X(_05588_));
 sky130_fd_sc_hd__nand2_1 _12780_ (.A(_05587_),
    .B(_05588_),
    .Y(_05589_));
 sky130_fd_sc_hd__xnor2_1 _12781_ (.A(_05547_),
    .B(_05589_),
    .Y(_05590_));
 sky130_fd_sc_hd__a21oi_2 _12782_ (.A1(_05562_),
    .A2(_05554_),
    .B1(_05590_),
    .Y(_05591_));
 sky130_fd_sc_hd__and3_1 _12783_ (.A(_05562_),
    .B(_05554_),
    .C(_05590_),
    .X(_05592_));
 sky130_fd_sc_hd__a211oi_2 _12784_ (.A1(_05556_),
    .A2(_05558_),
    .B1(_05591_),
    .C1(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__o211a_1 _12785_ (.A1(_05591_),
    .A2(_05592_),
    .B1(_05556_),
    .C1(_05558_),
    .X(_05594_));
 sky130_fd_sc_hd__or3_1 _12786_ (.A(_05327_),
    .B(_05593_),
    .C(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__a21oi_1 _12787_ (.A1(_05561_),
    .A2(_05595_),
    .B1(_05440_),
    .Y(_00313_));
 sky130_fd_sc_hd__a22o_1 _12788_ (.A1(_05304_),
    .A2(_05567_),
    .B1(_05297_),
    .B2(_05302_),
    .X(_05596_));
 sky130_fd_sc_hd__inv_2 _12789_ (.A(_05296_),
    .Y(_05597_));
 sky130_fd_sc_hd__or4_1 _12790_ (.A(_05447_),
    .B(_05449_),
    .C(_05292_),
    .D(_05597_),
    .X(_05598_));
 sky130_fd_sc_hd__nand2_1 _12791_ (.A(_05596_),
    .B(_05598_),
    .Y(_05599_));
 sky130_fd_sc_hd__nand2_1 _12792_ (.A(_05298_),
    .B(_05301_),
    .Y(_05600_));
 sky130_fd_sc_hd__xnor2_1 _12793_ (.A(_05599_),
    .B(_05600_),
    .Y(_05601_));
 sky130_fd_sc_hd__o21a_1 _12794_ (.A1(_05569_),
    .A2(_05570_),
    .B1(_05568_),
    .X(_05602_));
 sky130_fd_sc_hd__xor2_1 _12795_ (.A(_05601_),
    .B(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__o21ai_1 _12796_ (.A1(_05293_),
    .A2(_05288_),
    .B1(_05306_),
    .Y(_05604_));
 sky130_fd_sc_hd__and3_1 _12797_ (.A(_05293_),
    .B(_05288_),
    .C(_05305_),
    .X(_05605_));
 sky130_fd_sc_hd__nor3_1 _12798_ (.A(_05538_),
    .B(_05604_),
    .C(_05605_),
    .Y(_05606_));
 sky130_fd_sc_hd__o21a_1 _12799_ (.A1(_05604_),
    .A2(_05605_),
    .B1(_05538_),
    .X(_05607_));
 sky130_fd_sc_hd__nor2_2 _12800_ (.A(_05606_),
    .B(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__or2_1 _12801_ (.A(_05603_),
    .B(_05608_),
    .X(_05609_));
 sky130_fd_sc_hd__nand2_1 _12802_ (.A(_05603_),
    .B(_05608_),
    .Y(_05610_));
 sky130_fd_sc_hd__and2_1 _12803_ (.A(_05609_),
    .B(_05610_),
    .X(_05611_));
 sky130_fd_sc_hd__or2b_1 _12804_ (.A(_05573_),
    .B_N(_05577_),
    .X(_05612_));
 sky130_fd_sc_hd__o21a_1 _12805_ (.A1(_05571_),
    .A2(_05572_),
    .B1(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__xnor2_1 _12806_ (.A(_05611_),
    .B(_05613_),
    .Y(_05614_));
 sky130_fd_sc_hd__o21ba_1 _12807_ (.A1(_05538_),
    .A2(_05574_),
    .B1_N(_05575_),
    .X(_05615_));
 sky130_fd_sc_hd__nor2_1 _12808_ (.A(_05507_),
    .B(_05615_),
    .Y(_05616_));
 sky130_fd_sc_hd__and2_1 _12809_ (.A(_05507_),
    .B(_05615_),
    .X(_05617_));
 sky130_fd_sc_hd__nor2_1 _12810_ (.A(_05616_),
    .B(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__and2_1 _12811_ (.A(_05614_),
    .B(_05618_),
    .X(_05619_));
 sky130_fd_sc_hd__nor2_1 _12812_ (.A(_05614_),
    .B(_05618_),
    .Y(_05620_));
 sky130_fd_sc_hd__or2_1 _12813_ (.A(_05619_),
    .B(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__nand2_1 _12814_ (.A(_05579_),
    .B(_05585_),
    .Y(_05622_));
 sky130_fd_sc_hd__xor2_1 _12815_ (.A(_05621_),
    .B(_05622_),
    .X(_05623_));
 sky130_fd_sc_hd__or2_1 _12816_ (.A(_05582_),
    .B(_05623_),
    .X(_05624_));
 sky130_fd_sc_hd__nand2_1 _12817_ (.A(_05582_),
    .B(_05623_),
    .Y(_05625_));
 sky130_fd_sc_hd__nand2_1 _12818_ (.A(_05624_),
    .B(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__o21ai_1 _12819_ (.A1(_05547_),
    .A2(_05589_),
    .B1(_05587_),
    .Y(_05627_));
 sky130_fd_sc_hd__xnor2_1 _12820_ (.A(_05626_),
    .B(_05627_),
    .Y(_05628_));
 sky130_fd_sc_hd__o21ai_2 _12821_ (.A1(_05591_),
    .A2(_05593_),
    .B1(_05628_),
    .Y(_05629_));
 sky130_fd_sc_hd__or3_1 _12822_ (.A(_05591_),
    .B(_05593_),
    .C(_05628_),
    .X(_05630_));
 sky130_fd_sc_hd__a21o_1 _12823_ (.A1(_05629_),
    .A2(_05630_),
    .B1(_05328_),
    .X(_05631_));
 sky130_fd_sc_hd__o211a_1 _12824_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[11] ),
    .A2(_05314_),
    .B1(_05631_),
    .C1(_05308_),
    .X(_00314_));
 sky130_fd_sc_hd__clkbuf_8 _12825_ (.A(_04867_),
    .X(_05632_));
 sky130_fd_sc_hd__buf_8 _12826_ (.A(_05325_),
    .X(_05633_));
 sky130_fd_sc_hd__buf_6 _12827_ (.A(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__or2b_1 _12828_ (.A(_05626_),
    .B_N(_05627_),
    .X(_05635_));
 sky130_fd_sc_hd__or3b_1 _12829_ (.A(_05619_),
    .B(_05620_),
    .C_N(_05622_),
    .X(_05636_));
 sky130_fd_sc_hd__and2b_1 _12830_ (.A_N(_05613_),
    .B(_05611_),
    .X(_05637_));
 sky130_fd_sc_hd__or2_1 _12831_ (.A(_05601_),
    .B(_05602_),
    .X(_05638_));
 sky130_fd_sc_hd__a22o_1 _12832_ (.A1(_05304_),
    .A2(_05597_),
    .B1(_05301_),
    .B2(_05302_),
    .X(_05639_));
 sky130_fd_sc_hd__and2b_1 _12833_ (.A_N(_05267_),
    .B(\top_inst.skew_buff_inst.row[0].output_reg[6] ),
    .X(_05640_));
 sky130_fd_sc_hd__a21oi_2 _12834_ (.A1(\top_inst.axis_in_inst.inbuf_bus[6] ),
    .A2(_05267_),
    .B1(_05640_),
    .Y(_05641_));
 sky130_fd_sc_hd__or4_1 _12835_ (.A(_05447_),
    .B(_05449_),
    .C(_05297_),
    .D(_05641_),
    .X(_05642_));
 sky130_fd_sc_hd__nand2_1 _12836_ (.A(_05639_),
    .B(_05642_),
    .Y(_05643_));
 sky130_fd_sc_hd__nand2_2 _12837_ (.A(_05298_),
    .B(_05306_),
    .Y(_05644_));
 sky130_fd_sc_hd__xnor2_1 _12838_ (.A(_05643_),
    .B(_05644_),
    .Y(_05645_));
 sky130_fd_sc_hd__o21a_1 _12839_ (.A1(_05599_),
    .A2(_05600_),
    .B1(_05598_),
    .X(_05646_));
 sky130_fd_sc_hd__nor2_1 _12840_ (.A(_05645_),
    .B(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__and2_1 _12841_ (.A(_05645_),
    .B(_05646_),
    .X(_05648_));
 sky130_fd_sc_hd__nor2_1 _12842_ (.A(_05647_),
    .B(_05648_),
    .Y(_05649_));
 sky130_fd_sc_hd__xnor2_1 _12843_ (.A(_05608_),
    .B(_05649_),
    .Y(_05650_));
 sky130_fd_sc_hd__a21o_1 _12844_ (.A1(_05638_),
    .A2(_05610_),
    .B1(_05650_),
    .X(_05651_));
 sky130_fd_sc_hd__nand3_1 _12845_ (.A(_05638_),
    .B(_05610_),
    .C(_05650_),
    .Y(_05652_));
 sky130_fd_sc_hd__nand2_1 _12846_ (.A(_05651_),
    .B(_05652_),
    .Y(_05653_));
 sky130_fd_sc_hd__o21a_1 _12847_ (.A1(_05280_),
    .A2(_05273_),
    .B1(_05306_),
    .X(_05654_));
 sky130_fd_sc_hd__o21a_2 _12848_ (.A1(_05605_),
    .A2(_05606_),
    .B1(_05654_),
    .X(_05655_));
 sky130_fd_sc_hd__or3_1 _12849_ (.A(_05654_),
    .B(_05605_),
    .C(_05606_),
    .X(_05656_));
 sky130_fd_sc_hd__or2b_1 _12850_ (.A(_05655_),
    .B_N(_05656_),
    .X(_05657_));
 sky130_fd_sc_hd__clkbuf_2 _12851_ (.A(_05657_),
    .X(_05658_));
 sky130_fd_sc_hd__xor2_1 _12852_ (.A(_05653_),
    .B(_05658_),
    .X(_05659_));
 sky130_fd_sc_hd__o21ai_1 _12853_ (.A1(_05637_),
    .A2(_05619_),
    .B1(_05659_),
    .Y(_05660_));
 sky130_fd_sc_hd__or3_1 _12854_ (.A(_05637_),
    .B(_05619_),
    .C(_05659_),
    .X(_05661_));
 sky130_fd_sc_hd__and2_1 _12855_ (.A(_05660_),
    .B(_05661_),
    .X(_05662_));
 sky130_fd_sc_hd__xnor2_1 _12856_ (.A(_05616_),
    .B(_05662_),
    .Y(_05663_));
 sky130_fd_sc_hd__a21oi_1 _12857_ (.A1(_05636_),
    .A2(_05624_),
    .B1(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__and3_1 _12858_ (.A(_05636_),
    .B(_05624_),
    .C(_05663_),
    .X(_05665_));
 sky130_fd_sc_hd__or2_1 _12859_ (.A(_05664_),
    .B(_05665_),
    .X(_05666_));
 sky130_fd_sc_hd__a21oi_2 _12860_ (.A1(_05635_),
    .A2(_05629_),
    .B1(_05666_),
    .Y(_05667_));
 sky130_fd_sc_hd__a31o_1 _12861_ (.A1(_05635_),
    .A2(_05629_),
    .A3(_05666_),
    .B1(_05633_),
    .X(_05668_));
 sky130_fd_sc_hd__o2bb2a_1 _12862_ (.A1_N(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[12] ),
    .A2_N(_05634_),
    .B1(_05667_),
    .B2(_05668_),
    .X(_05669_));
 sky130_fd_sc_hd__nor2_1 _12863_ (.A(_05632_),
    .B(_05669_),
    .Y(_00315_));
 sky130_fd_sc_hd__nand2_1 _12864_ (.A(_05616_),
    .B(_05662_),
    .Y(_05670_));
 sky130_fd_sc_hd__or2_1 _12865_ (.A(_05643_),
    .B(_05644_),
    .X(_05671_));
 sky130_fd_sc_hd__and2_1 _12866_ (.A(_05302_),
    .B(_05305_),
    .X(_05672_));
 sky130_fd_sc_hd__a21oi_1 _12867_ (.A1(_05304_),
    .A2(_05641_),
    .B1(_05672_),
    .Y(_05673_));
 sky130_fd_sc_hd__and3_1 _12868_ (.A(_05304_),
    .B(_05641_),
    .C(_05672_),
    .X(_05674_));
 sky130_fd_sc_hd__or2_1 _12869_ (.A(_05673_),
    .B(_05674_),
    .X(_05675_));
 sky130_fd_sc_hd__xnor2_1 _12870_ (.A(_05644_),
    .B(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__a21o_1 _12871_ (.A1(_05642_),
    .A2(_05671_),
    .B1(_05676_),
    .X(_05677_));
 sky130_fd_sc_hd__nand3_1 _12872_ (.A(_05642_),
    .B(_05671_),
    .C(_05676_),
    .Y(_05678_));
 sky130_fd_sc_hd__and2_1 _12873_ (.A(_05677_),
    .B(_05678_),
    .X(_05679_));
 sky130_fd_sc_hd__nand2_1 _12874_ (.A(_05608_),
    .B(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hd__or2_1 _12875_ (.A(_05608_),
    .B(_05679_),
    .X(_05681_));
 sky130_fd_sc_hd__nand2_1 _12876_ (.A(_05680_),
    .B(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__a21o_1 _12877_ (.A1(_05608_),
    .A2(_05649_),
    .B1(_05647_),
    .X(_05683_));
 sky130_fd_sc_hd__xor2_1 _12878_ (.A(_05682_),
    .B(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__xnor2_1 _12879_ (.A(_05658_),
    .B(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__o21a_1 _12880_ (.A1(_05653_),
    .A2(_05658_),
    .B1(_05651_),
    .X(_05686_));
 sky130_fd_sc_hd__nor2_1 _12881_ (.A(_05685_),
    .B(_05686_),
    .Y(_05687_));
 sky130_fd_sc_hd__and2_1 _12882_ (.A(_05685_),
    .B(_05686_),
    .X(_05688_));
 sky130_fd_sc_hd__nor2_1 _12883_ (.A(_05687_),
    .B(_05688_),
    .Y(_05689_));
 sky130_fd_sc_hd__xnor2_1 _12884_ (.A(_05655_),
    .B(_05689_),
    .Y(_05690_));
 sky130_fd_sc_hd__a21o_1 _12885_ (.A1(_05660_),
    .A2(_05670_),
    .B1(_05690_),
    .X(_05691_));
 sky130_fd_sc_hd__nand3_1 _12886_ (.A(_05660_),
    .B(_05670_),
    .C(_05690_),
    .Y(_05692_));
 sky130_fd_sc_hd__and2_1 _12887_ (.A(_05691_),
    .B(_05692_),
    .X(_05693_));
 sky130_fd_sc_hd__or3_1 _12888_ (.A(_05664_),
    .B(_05667_),
    .C(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__o21ai_1 _12889_ (.A1(_05664_),
    .A2(_05667_),
    .B1(_05693_),
    .Y(_05695_));
 sky130_fd_sc_hd__and2_1 _12890_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[13] ),
    .B(_05326_),
    .X(_05696_));
 sky130_fd_sc_hd__a31o_1 _12891_ (.A1(_05335_),
    .A2(_05694_),
    .A3(_05695_),
    .B1(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__and2_1 _12892_ (.A(_05352_),
    .B(_05697_),
    .X(_05698_));
 sky130_fd_sc_hd__clkbuf_1 _12893_ (.A(_05698_),
    .X(_00316_));
 sky130_fd_sc_hd__nand2_1 _12894_ (.A(net998),
    .B(_05403_),
    .Y(_05699_));
 sky130_fd_sc_hd__nand2_1 _12895_ (.A(_05302_),
    .B(_05306_),
    .Y(_05700_));
 sky130_fd_sc_hd__o211a_1 _12896_ (.A1(_05447_),
    .A2(_05306_),
    .B1(_05644_),
    .C1(_05700_),
    .X(_05701_));
 sky130_fd_sc_hd__o21ba_1 _12897_ (.A1(_05644_),
    .A2(_05673_),
    .B1_N(_05674_),
    .X(_05702_));
 sky130_fd_sc_hd__a21oi_1 _12898_ (.A1(_05298_),
    .A2(_05672_),
    .B1(_05702_),
    .Y(_05703_));
 sky130_fd_sc_hd__nor2_1 _12899_ (.A(_05701_),
    .B(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hd__xnor2_1 _12900_ (.A(_05608_),
    .B(_05704_),
    .Y(_05705_));
 sky130_fd_sc_hd__a21o_1 _12901_ (.A1(_05677_),
    .A2(_05680_),
    .B1(_05705_),
    .X(_05706_));
 sky130_fd_sc_hd__nand3_1 _12902_ (.A(_05677_),
    .B(_05680_),
    .C(_05705_),
    .Y(_05707_));
 sky130_fd_sc_hd__and2_1 _12903_ (.A(_05706_),
    .B(_05707_),
    .X(_05708_));
 sky130_fd_sc_hd__xor2_1 _12904_ (.A(_05658_),
    .B(_05708_),
    .X(_05709_));
 sky130_fd_sc_hd__or2b_1 _12905_ (.A(_05682_),
    .B_N(_05683_),
    .X(_05710_));
 sky130_fd_sc_hd__o21ai_1 _12906_ (.A1(_05658_),
    .A2(_05684_),
    .B1(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__xnor2_1 _12907_ (.A(_05709_),
    .B(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__xnor2_1 _12908_ (.A(_05655_),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__a21oi_1 _12909_ (.A1(_05655_),
    .A2(_05689_),
    .B1(_05687_),
    .Y(_05714_));
 sky130_fd_sc_hd__or2_1 _12910_ (.A(_05713_),
    .B(_05714_),
    .X(_05715_));
 sky130_fd_sc_hd__nand2_1 _12911_ (.A(_05713_),
    .B(_05714_),
    .Y(_05716_));
 sky130_fd_sc_hd__nand2_1 _12912_ (.A(_05715_),
    .B(_05716_),
    .Y(_05717_));
 sky130_fd_sc_hd__and3_1 _12913_ (.A(_05691_),
    .B(_05695_),
    .C(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__a21o_1 _12914_ (.A1(_05691_),
    .A2(_05695_),
    .B1(_05717_),
    .X(_05719_));
 sky130_fd_sc_hd__or3b_1 _12915_ (.A(_05718_),
    .B(_05406_),
    .C_N(_05719_),
    .X(_05720_));
 sky130_fd_sc_hd__a21oi_1 _12916_ (.A1(_05699_),
    .A2(_05720_),
    .B1(_05440_),
    .Y(_00317_));
 sky130_fd_sc_hd__and2b_1 _12917_ (.A_N(_05709_),
    .B(_05711_),
    .X(_05721_));
 sky130_fd_sc_hd__a21o_1 _12918_ (.A1(_05655_),
    .A2(_05712_),
    .B1(_05721_),
    .X(_05722_));
 sky130_fd_sc_hd__mux2_1 _12919_ (.A0(_05703_),
    .A1(_05701_),
    .S(_05608_),
    .X(_05723_));
 sky130_fd_sc_hd__xnor2_1 _12920_ (.A(_05722_),
    .B(_05723_),
    .Y(_05724_));
 sky130_fd_sc_hd__inv_2 _12921_ (.A(_05708_),
    .Y(_05725_));
 sky130_fd_sc_hd__o21ai_1 _12922_ (.A1(_05658_),
    .A2(_05725_),
    .B1(_05656_),
    .Y(_05726_));
 sky130_fd_sc_hd__mux2_1 _12923_ (.A0(_05656_),
    .A1(_05726_),
    .S(_05706_),
    .X(_05727_));
 sky130_fd_sc_hd__xor2_1 _12924_ (.A(_05701_),
    .B(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__xnor2_1 _12925_ (.A(_05724_),
    .B(_05728_),
    .Y(_05729_));
 sky130_fd_sc_hd__clkbuf_8 _12926_ (.A(_05324_),
    .X(_05730_));
 sky130_fd_sc_hd__buf_6 _12927_ (.A(_05730_),
    .X(_05731_));
 sky130_fd_sc_hd__buf_12 _12928_ (.A(_05731_),
    .X(_05732_));
 sky130_fd_sc_hd__a31o_1 _12929_ (.A1(_05715_),
    .A2(_05719_),
    .A3(_05729_),
    .B1(_05732_),
    .X(_05733_));
 sky130_fd_sc_hd__o211a_1 _12930_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[15] ),
    .A2(_05314_),
    .B1(_05733_),
    .C1(_05308_),
    .X(_00318_));
 sky130_fd_sc_hd__buf_4 _12931_ (.A(\top_inst.grid_inst.data_path_wires[1][0] ),
    .X(_05734_));
 sky130_fd_sc_hd__clkbuf_4 _12932_ (.A(_04865_),
    .X(_05735_));
 sky130_fd_sc_hd__clkbuf_8 _12933_ (.A(_04858_),
    .X(_05736_));
 sky130_fd_sc_hd__or2_1 _12934_ (.A(_05736_),
    .B(_05272_),
    .X(_05737_));
 sky130_fd_sc_hd__o211a_1 _12935_ (.A1(_05734_),
    .A2(_05735_),
    .B1(_05737_),
    .C1(_05308_),
    .X(_00319_));
 sky130_fd_sc_hd__clkbuf_4 _12936_ (.A(\top_inst.grid_inst.data_path_wires[1][1] ),
    .X(_05738_));
 sky130_fd_sc_hd__buf_6 _12937_ (.A(_04864_),
    .X(_05739_));
 sky130_fd_sc_hd__nand2_1 _12938_ (.A(_05739_),
    .B(_05488_),
    .Y(_05740_));
 sky130_fd_sc_hd__o211a_1 _12939_ (.A1(_05738_),
    .A2(_05735_),
    .B1(_05740_),
    .C1(_05308_),
    .X(_00320_));
 sky130_fd_sc_hd__clkbuf_4 _12940_ (.A(\top_inst.grid_inst.data_path_wires[1][2] ),
    .X(_05741_));
 sky130_fd_sc_hd__nand2_1 _12941_ (.A(_05739_),
    .B(_05490_),
    .Y(_05742_));
 sky130_fd_sc_hd__clkbuf_4 _12942_ (.A(_05260_),
    .X(_05743_));
 sky130_fd_sc_hd__o211a_1 _12943_ (.A1(_05741_),
    .A2(_05735_),
    .B1(_05742_),
    .C1(_05743_),
    .X(_00321_));
 sky130_fd_sc_hd__buf_4 _12944_ (.A(\top_inst.grid_inst.data_path_wires[1][3] ),
    .X(_05744_));
 sky130_fd_sc_hd__nand2_1 _12945_ (.A(_05739_),
    .B(_05528_),
    .Y(_05745_));
 sky130_fd_sc_hd__o211a_1 _12946_ (.A1(_05744_),
    .A2(_05735_),
    .B1(_05745_),
    .C1(_05743_),
    .X(_00322_));
 sky130_fd_sc_hd__clkbuf_4 _12947_ (.A(\top_inst.grid_inst.data_path_wires[1][4] ),
    .X(_05746_));
 sky130_fd_sc_hd__nand2_1 _12948_ (.A(_05739_),
    .B(_05567_),
    .Y(_05747_));
 sky130_fd_sc_hd__o211a_1 _12949_ (.A1(_05746_),
    .A2(_05735_),
    .B1(_05747_),
    .C1(_05743_),
    .X(_00323_));
 sky130_fd_sc_hd__clkbuf_4 _12950_ (.A(\top_inst.grid_inst.data_path_wires[1][5] ),
    .X(_05748_));
 sky130_fd_sc_hd__nand2_1 _12951_ (.A(_05739_),
    .B(_05597_),
    .Y(_05749_));
 sky130_fd_sc_hd__o211a_1 _12952_ (.A1(_05748_),
    .A2(_05735_),
    .B1(_05749_),
    .C1(_05743_),
    .X(_00324_));
 sky130_fd_sc_hd__buf_2 _12953_ (.A(\top_inst.grid_inst.data_path_wires[1][6] ),
    .X(_05750_));
 sky130_fd_sc_hd__clkbuf_4 _12954_ (.A(_05750_),
    .X(_05751_));
 sky130_fd_sc_hd__nand2_1 _12955_ (.A(_05739_),
    .B(_05641_),
    .Y(_05752_));
 sky130_fd_sc_hd__o211a_1 _12956_ (.A1(_05751_),
    .A2(_05735_),
    .B1(_05752_),
    .C1(_05743_),
    .X(_00325_));
 sky130_fd_sc_hd__clkbuf_4 _12957_ (.A(\top_inst.grid_inst.data_path_wires[1][7] ),
    .X(_05753_));
 sky130_fd_sc_hd__or2_1 _12958_ (.A(_05736_),
    .B(_05306_),
    .X(_05754_));
 sky130_fd_sc_hd__o211a_1 _12959_ (.A1(_05753_),
    .A2(_05735_),
    .B1(_05754_),
    .C1(_05743_),
    .X(_00326_));
 sky130_fd_sc_hd__clkbuf_8 _12960_ (.A(_05268_),
    .X(_05755_));
 sky130_fd_sc_hd__clkbuf_4 _12961_ (.A(_05755_),
    .X(_05756_));
 sky130_fd_sc_hd__clkbuf_4 _12962_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[0] ),
    .X(_05757_));
 sky130_fd_sc_hd__or2_1 _12963_ (.A(_05757_),
    .B(_05294_),
    .X(_05758_));
 sky130_fd_sc_hd__o211a_1 _12964_ (.A1(_05734_),
    .A2(_05756_),
    .B1(_05758_),
    .C1(_05743_),
    .X(_00327_));
 sky130_fd_sc_hd__clkbuf_4 _12965_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[1] ),
    .X(_05759_));
 sky130_fd_sc_hd__or2_1 _12966_ (.A(_05759_),
    .B(_05294_),
    .X(_05760_));
 sky130_fd_sc_hd__o211a_1 _12967_ (.A1(_05738_),
    .A2(_05756_),
    .B1(_05760_),
    .C1(_05743_),
    .X(_00328_));
 sky130_fd_sc_hd__clkbuf_4 _12968_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[2] ),
    .X(_05761_));
 sky130_fd_sc_hd__or2_1 _12969_ (.A(_05761_),
    .B(_05294_),
    .X(_05762_));
 sky130_fd_sc_hd__o211a_1 _12970_ (.A1(_05741_),
    .A2(_05756_),
    .B1(_05762_),
    .C1(_05743_),
    .X(_00329_));
 sky130_fd_sc_hd__clkbuf_4 _12971_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[3] ),
    .X(_05763_));
 sky130_fd_sc_hd__or2_1 _12972_ (.A(_05763_),
    .B(_05294_),
    .X(_05764_));
 sky130_fd_sc_hd__o211a_1 _12973_ (.A1(_05744_),
    .A2(_05756_),
    .B1(_05764_),
    .C1(_05743_),
    .X(_00330_));
 sky130_fd_sc_hd__clkbuf_4 _12974_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[4] ),
    .X(_05765_));
 sky130_fd_sc_hd__or2_1 _12975_ (.A(_05765_),
    .B(_05294_),
    .X(_05766_));
 sky130_fd_sc_hd__clkbuf_4 _12976_ (.A(_05260_),
    .X(_05767_));
 sky130_fd_sc_hd__o211a_1 _12977_ (.A1(_05746_),
    .A2(_05756_),
    .B1(_05766_),
    .C1(_05767_),
    .X(_00331_));
 sky130_fd_sc_hd__clkbuf_4 _12978_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[5] ),
    .X(_05768_));
 sky130_fd_sc_hd__or2_1 _12979_ (.A(_05768_),
    .B(_05294_),
    .X(_05769_));
 sky130_fd_sc_hd__o211a_1 _12980_ (.A1(_05748_),
    .A2(_05756_),
    .B1(_05769_),
    .C1(_05767_),
    .X(_00332_));
 sky130_fd_sc_hd__buf_2 _12981_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[6] ),
    .X(_05770_));
 sky130_fd_sc_hd__or2_1 _12982_ (.A(_05770_),
    .B(_05294_),
    .X(_05771_));
 sky130_fd_sc_hd__o211a_1 _12983_ (.A1(_05751_),
    .A2(_05756_),
    .B1(_05771_),
    .C1(_05767_),
    .X(_00333_));
 sky130_fd_sc_hd__buf_4 _12984_ (.A(_05274_),
    .X(_05772_));
 sky130_fd_sc_hd__clkbuf_4 _12985_ (.A(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__or2_1 _12986_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[7] ),
    .B(_05773_),
    .X(_05774_));
 sky130_fd_sc_hd__o211a_1 _12987_ (.A1(_05753_),
    .A2(_05756_),
    .B1(_05774_),
    .C1(_05767_),
    .X(_00334_));
 sky130_fd_sc_hd__nand2_1 _12988_ (.A(_05734_),
    .B(_05757_),
    .Y(_05775_));
 sky130_fd_sc_hd__nand2_1 _12989_ (.A(_05317_),
    .B(_05775_),
    .Y(_05776_));
 sky130_fd_sc_hd__o211a_1 _12990_ (.A1(net1044),
    .A2(_05314_),
    .B1(_05776_),
    .C1(_05767_),
    .X(_00335_));
 sky130_fd_sc_hd__nand2_1 _12991_ (.A(_05738_),
    .B(_05759_),
    .Y(_05777_));
 sky130_fd_sc_hd__a22o_1 _12992_ (.A1(_05734_),
    .A2(_05759_),
    .B1(_05757_),
    .B2(_05738_),
    .X(_05778_));
 sky130_fd_sc_hd__o21ai_1 _12993_ (.A1(_05775_),
    .A2(_05777_),
    .B1(_05778_),
    .Y(_05779_));
 sky130_fd_sc_hd__nand2_1 _12994_ (.A(_05317_),
    .B(_05779_),
    .Y(_05780_));
 sky130_fd_sc_hd__o211a_1 _12995_ (.A1(net1060),
    .A2(_05314_),
    .B1(_05780_),
    .C1(_05767_),
    .X(_00336_));
 sky130_fd_sc_hd__nand2_1 _12996_ (.A(_05741_),
    .B(_05757_),
    .Y(_05781_));
 sky130_fd_sc_hd__and3_1 _12997_ (.A(_05738_),
    .B(_05759_),
    .C(_05775_),
    .X(_05782_));
 sky130_fd_sc_hd__xnor2_1 _12998_ (.A(_05781_),
    .B(_05782_),
    .Y(_05783_));
 sky130_fd_sc_hd__a21oi_1 _12999_ (.A1(_05734_),
    .A2(_05761_),
    .B1(_05783_),
    .Y(_05784_));
 sky130_fd_sc_hd__and3_1 _13000_ (.A(_05734_),
    .B(_05761_),
    .C(_05783_),
    .X(_05785_));
 sky130_fd_sc_hd__o21ai_1 _13001_ (.A1(_05784_),
    .A2(_05785_),
    .B1(_05336_),
    .Y(_05786_));
 sky130_fd_sc_hd__o211a_1 _13002_ (.A1(net1087),
    .A2(_05314_),
    .B1(_05786_),
    .C1(_05767_),
    .X(_00337_));
 sky130_fd_sc_hd__buf_8 _13003_ (.A(_05312_),
    .X(_05787_));
 sky130_fd_sc_hd__buf_4 _13004_ (.A(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__a22oi_1 _13005_ (.A1(_05734_),
    .A2(_05763_),
    .B1(_05761_),
    .B2(_05738_),
    .Y(_05789_));
 sky130_fd_sc_hd__and4_1 _13006_ (.A(\top_inst.grid_inst.data_path_wires[1][1] ),
    .B(\top_inst.grid_inst.data_path_wires[1][0] ),
    .C(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[3] ),
    .D(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[2] ),
    .X(_05790_));
 sky130_fd_sc_hd__or2_1 _13007_ (.A(_05789_),
    .B(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__and4_1 _13008_ (.A(\top_inst.grid_inst.data_path_wires[1][3] ),
    .B(\top_inst.grid_inst.data_path_wires[1][2] ),
    .C(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[0] ),
    .X(_05792_));
 sky130_fd_sc_hd__o21a_1 _13009_ (.A1(_05777_),
    .A2(_05781_),
    .B1(_05792_),
    .X(_05793_));
 sky130_fd_sc_hd__a22o_1 _13010_ (.A1(_05741_),
    .A2(_05759_),
    .B1(_05757_),
    .B2(_05744_),
    .X(_05794_));
 sky130_fd_sc_hd__or3_1 _13011_ (.A(_05777_),
    .B(_05781_),
    .C(_05792_),
    .X(_05795_));
 sky130_fd_sc_hd__and3b_1 _13012_ (.A_N(_05793_),
    .B(_05794_),
    .C(_05795_),
    .X(_05796_));
 sky130_fd_sc_hd__xnor2_1 _13013_ (.A(_05791_),
    .B(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__nor3_1 _13014_ (.A(_05741_),
    .B(_05775_),
    .C(_05777_),
    .Y(_05798_));
 sky130_fd_sc_hd__nor3_1 _13015_ (.A(_05785_),
    .B(_05797_),
    .C(_05798_),
    .Y(_05799_));
 sky130_fd_sc_hd__o21a_1 _13016_ (.A1(_05785_),
    .A2(_05798_),
    .B1(_05797_),
    .X(_05800_));
 sky130_fd_sc_hd__o21ai_1 _13017_ (.A1(_05799_),
    .A2(_05800_),
    .B1(_05336_),
    .Y(_05801_));
 sky130_fd_sc_hd__o211a_1 _13018_ (.A1(net1073),
    .A2(_05788_),
    .B1(_05801_),
    .C1(_05767_),
    .X(_00338_));
 sky130_fd_sc_hd__and2b_1 _13019_ (.A_N(_05791_),
    .B(_05796_),
    .X(_05802_));
 sky130_fd_sc_hd__inv_2 _13020_ (.A(_05792_),
    .Y(_05803_));
 sky130_fd_sc_hd__nand4_1 _13021_ (.A(\top_inst.grid_inst.data_path_wires[1][4] ),
    .B(\top_inst.grid_inst.data_path_wires[1][3] ),
    .C(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[0] ),
    .Y(_05804_));
 sky130_fd_sc_hd__a22o_1 _13022_ (.A1(\top_inst.grid_inst.data_path_wires[1][3] ),
    .A2(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[1][4] ),
    .X(_05805_));
 sky130_fd_sc_hd__and3_1 _13023_ (.A(_05790_),
    .B(_05804_),
    .C(_05805_),
    .X(_05806_));
 sky130_fd_sc_hd__a21oi_1 _13024_ (.A1(_05804_),
    .A2(_05805_),
    .B1(_05790_),
    .Y(_05807_));
 sky130_fd_sc_hd__nor2_1 _13025_ (.A(_05806_),
    .B(_05807_),
    .Y(_05808_));
 sky130_fd_sc_hd__xnor2_1 _13026_ (.A(_05803_),
    .B(_05808_),
    .Y(_05809_));
 sky130_fd_sc_hd__nand2_1 _13027_ (.A(_05741_),
    .B(_05761_),
    .Y(_05810_));
 sky130_fd_sc_hd__and3_1 _13028_ (.A(\top_inst.grid_inst.data_path_wires[1][1] ),
    .B(\top_inst.grid_inst.data_path_wires[1][0] ),
    .C(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[3] ),
    .X(_05811_));
 sky130_fd_sc_hd__a22o_1 _13029_ (.A1(\top_inst.grid_inst.data_path_wires[1][0] ),
    .A2(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[1][1] ),
    .X(_05812_));
 sky130_fd_sc_hd__a21bo_1 _13030_ (.A1(_05765_),
    .A2(_05811_),
    .B1_N(_05812_),
    .X(_05813_));
 sky130_fd_sc_hd__xor2_1 _13031_ (.A(_05810_),
    .B(_05813_),
    .X(_05814_));
 sky130_fd_sc_hd__xor2_1 _13032_ (.A(_05809_),
    .B(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__xnor2_1 _13033_ (.A(_05802_),
    .B(_05815_),
    .Y(_05816_));
 sky130_fd_sc_hd__xor2_1 _13034_ (.A(_05795_),
    .B(_05816_),
    .X(_05817_));
 sky130_fd_sc_hd__nand2_1 _13035_ (.A(_05800_),
    .B(_05817_),
    .Y(_05818_));
 sky130_fd_sc_hd__o21a_1 _13036_ (.A1(_05800_),
    .A2(_05817_),
    .B1(_05315_),
    .X(_05819_));
 sky130_fd_sc_hd__a22o_1 _13037_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[4] ),
    .A2(_05354_),
    .B1(_05818_),
    .B2(_05819_),
    .X(_05820_));
 sky130_fd_sc_hd__and2_1 _13038_ (.A(_05352_),
    .B(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__clkbuf_1 _13039_ (.A(_05821_),
    .X(_00339_));
 sky130_fd_sc_hd__and2_1 _13040_ (.A(_05809_),
    .B(_05814_),
    .X(_05822_));
 sky130_fd_sc_hd__nand2_1 _13041_ (.A(_05734_),
    .B(_05768_),
    .Y(_05823_));
 sky130_fd_sc_hd__a22o_1 _13042_ (.A1(\top_inst.grid_inst.data_path_wires[1][1] ),
    .A2(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[1][2] ),
    .X(_05824_));
 sky130_fd_sc_hd__nand4_1 _13043_ (.A(\top_inst.grid_inst.data_path_wires[1][2] ),
    .B(_05738_),
    .C(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[3] ),
    .Y(_05825_));
 sky130_fd_sc_hd__nand2_1 _13044_ (.A(_05824_),
    .B(_05825_),
    .Y(_05826_));
 sky130_fd_sc_hd__and2_1 _13045_ (.A(\top_inst.grid_inst.data_path_wires[1][3] ),
    .B(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[2] ),
    .X(_05827_));
 sky130_fd_sc_hd__xor2_2 _13046_ (.A(_05826_),
    .B(_05827_),
    .X(_05828_));
 sky130_fd_sc_hd__xor2_2 _13047_ (.A(_05823_),
    .B(_05828_),
    .X(_05829_));
 sky130_fd_sc_hd__and4_1 _13048_ (.A(_05746_),
    .B(_05744_),
    .C(_05759_),
    .D(_05757_),
    .X(_05830_));
 sky130_fd_sc_hd__a32o_1 _13049_ (.A1(\top_inst.grid_inst.data_path_wires[1][2] ),
    .A2(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[2] ),
    .A3(_05812_),
    .B1(_05811_),
    .B2(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[4] ),
    .X(_05831_));
 sky130_fd_sc_hd__and4_1 _13050_ (.A(\top_inst.grid_inst.data_path_wires[1][5] ),
    .B(\top_inst.grid_inst.data_path_wires[1][4] ),
    .C(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[0] ),
    .X(_05832_));
 sky130_fd_sc_hd__a22oi_1 _13051_ (.A1(\top_inst.grid_inst.data_path_wires[1][4] ),
    .A2(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[1][5] ),
    .Y(_05833_));
 sky130_fd_sc_hd__nor2_1 _13052_ (.A(_05832_),
    .B(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__xor2_2 _13053_ (.A(_05831_),
    .B(_05834_),
    .X(_05835_));
 sky130_fd_sc_hd__xnor2_2 _13054_ (.A(_05830_),
    .B(_05835_),
    .Y(_05836_));
 sky130_fd_sc_hd__xor2_2 _13055_ (.A(_05829_),
    .B(_05836_),
    .X(_05837_));
 sky130_fd_sc_hd__xnor2_1 _13056_ (.A(_05822_),
    .B(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__o21ba_1 _13057_ (.A1(_05803_),
    .A2(_05807_),
    .B1_N(_05806_),
    .X(_05839_));
 sky130_fd_sc_hd__xor2_1 _13058_ (.A(_05838_),
    .B(_05839_),
    .X(_05840_));
 sky130_fd_sc_hd__nand2_1 _13059_ (.A(_05802_),
    .B(_05815_),
    .Y(_05841_));
 sky130_fd_sc_hd__o21a_1 _13060_ (.A1(_05795_),
    .A2(_05816_),
    .B1(_05841_),
    .X(_05842_));
 sky130_fd_sc_hd__xnor2_1 _13061_ (.A(_05840_),
    .B(_05842_),
    .Y(_05843_));
 sky130_fd_sc_hd__or2_1 _13062_ (.A(_05818_),
    .B(_05843_),
    .X(_05844_));
 sky130_fd_sc_hd__a21oi_1 _13063_ (.A1(_05818_),
    .A2(_05843_),
    .B1(_05399_),
    .Y(_05845_));
 sky130_fd_sc_hd__a22o_1 _13064_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[5] ),
    .A2(_05354_),
    .B1(_05844_),
    .B2(_05845_),
    .X(_05846_));
 sky130_fd_sc_hd__and2_1 _13065_ (.A(_05352_),
    .B(_05846_),
    .X(_05847_));
 sky130_fd_sc_hd__clkbuf_1 _13066_ (.A(_05847_),
    .X(_00340_));
 sky130_fd_sc_hd__or2_1 _13067_ (.A(_05840_),
    .B(_05842_),
    .X(_05848_));
 sky130_fd_sc_hd__nand2_1 _13068_ (.A(_05831_),
    .B(_05834_),
    .Y(_05849_));
 sky130_fd_sc_hd__nand2_1 _13069_ (.A(_05830_),
    .B(_05835_),
    .Y(_05850_));
 sky130_fd_sc_hd__inv_2 _13070_ (.A(_05829_),
    .Y(_05851_));
 sky130_fd_sc_hd__nor2_1 _13071_ (.A(_05851_),
    .B(_05836_),
    .Y(_05852_));
 sky130_fd_sc_hd__or2_1 _13072_ (.A(_05823_),
    .B(_05828_),
    .X(_05853_));
 sky130_fd_sc_hd__a22o_1 _13073_ (.A1(_05734_),
    .A2(_05770_),
    .B1(_05768_),
    .B2(_05738_),
    .X(_05854_));
 sky130_fd_sc_hd__nand4_2 _13074_ (.A(_05738_),
    .B(\top_inst.grid_inst.data_path_wires[1][0] ),
    .C(_05770_),
    .D(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[5] ),
    .Y(_05855_));
 sky130_fd_sc_hd__nand2_1 _13075_ (.A(_05854_),
    .B(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__a22o_1 _13076_ (.A1(\top_inst.grid_inst.data_path_wires[1][2] ),
    .A2(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[1][3] ),
    .X(_05857_));
 sky130_fd_sc_hd__nand4_2 _13077_ (.A(\top_inst.grid_inst.data_path_wires[1][3] ),
    .B(_05741_),
    .C(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[3] ),
    .Y(_05858_));
 sky130_fd_sc_hd__a22o_1 _13078_ (.A1(_05746_),
    .A2(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[2] ),
    .B1(_05857_),
    .B2(_05858_),
    .X(_05859_));
 sky130_fd_sc_hd__nand4_1 _13079_ (.A(_05746_),
    .B(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[2] ),
    .C(_05857_),
    .D(_05858_),
    .Y(_05860_));
 sky130_fd_sc_hd__nand2_1 _13080_ (.A(_05859_),
    .B(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__xnor2_2 _13081_ (.A(_05856_),
    .B(_05861_),
    .Y(_05862_));
 sky130_fd_sc_hd__xnor2_2 _13082_ (.A(_05853_),
    .B(_05862_),
    .Y(_05863_));
 sky130_fd_sc_hd__a21bo_1 _13083_ (.A1(_05824_),
    .A2(_05827_),
    .B1_N(_05825_),
    .X(_05864_));
 sky130_fd_sc_hd__and4_1 _13084_ (.A(_05750_),
    .B(\top_inst.grid_inst.data_path_wires[1][5] ),
    .C(_05759_),
    .D(_05757_),
    .X(_05865_));
 sky130_fd_sc_hd__a22oi_1 _13085_ (.A1(\top_inst.grid_inst.data_path_wires[1][5] ),
    .A2(_05759_),
    .B1(_05757_),
    .B2(_05750_),
    .Y(_05866_));
 sky130_fd_sc_hd__nor2_1 _13086_ (.A(_05865_),
    .B(_05866_),
    .Y(_05867_));
 sky130_fd_sc_hd__and2_1 _13087_ (.A(_05864_),
    .B(_05867_),
    .X(_05868_));
 sky130_fd_sc_hd__nor2_1 _13088_ (.A(_05864_),
    .B(_05867_),
    .Y(_05869_));
 sky130_fd_sc_hd__nor2_1 _13089_ (.A(_05868_),
    .B(_05869_),
    .Y(_05870_));
 sky130_fd_sc_hd__xnor2_2 _13090_ (.A(_05832_),
    .B(_05870_),
    .Y(_05871_));
 sky130_fd_sc_hd__xnor2_2 _13091_ (.A(_05863_),
    .B(_05871_),
    .Y(_05872_));
 sky130_fd_sc_hd__xor2_1 _13092_ (.A(_05852_),
    .B(_05872_),
    .X(_05873_));
 sky130_fd_sc_hd__a21oi_1 _13093_ (.A1(_05849_),
    .A2(_05850_),
    .B1(_05873_),
    .Y(_05874_));
 sky130_fd_sc_hd__and3_1 _13094_ (.A(_05849_),
    .B(_05850_),
    .C(_05873_),
    .X(_05875_));
 sky130_fd_sc_hd__inv_2 _13095_ (.A(_05837_),
    .Y(_05876_));
 sky130_fd_sc_hd__and2b_1 _13096_ (.A_N(_05839_),
    .B(_05838_),
    .X(_05877_));
 sky130_fd_sc_hd__a21oi_1 _13097_ (.A1(_05822_),
    .A2(_05876_),
    .B1(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__nor3_1 _13098_ (.A(_05874_),
    .B(_05875_),
    .C(_05878_),
    .Y(_05879_));
 sky130_fd_sc_hd__o21a_1 _13099_ (.A1(_05874_),
    .A2(_05875_),
    .B1(_05878_),
    .X(_05880_));
 sky130_fd_sc_hd__a211oi_2 _13100_ (.A1(_05848_),
    .A2(_05844_),
    .B1(net169),
    .C1(_05880_),
    .Y(_05881_));
 sky130_fd_sc_hd__o211a_1 _13101_ (.A1(net169),
    .A2(_05880_),
    .B1(_05848_),
    .C1(_05844_),
    .X(_05882_));
 sky130_fd_sc_hd__or2_1 _13102_ (.A(_05325_),
    .B(_05882_),
    .X(_05883_));
 sky130_fd_sc_hd__a2bb2o_1 _13103_ (.A1_N(_05881_),
    .A2_N(_05883_),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[6] ),
    .B2(_05327_),
    .X(_05884_));
 sky130_fd_sc_hd__and2_1 _13104_ (.A(_05352_),
    .B(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__clkbuf_1 _13105_ (.A(_05885_),
    .X(_00341_));
 sky130_fd_sc_hd__clkbuf_4 _13106_ (.A(_04869_),
    .X(_05886_));
 sky130_fd_sc_hd__buf_8 _13107_ (.A(_05315_),
    .X(_05887_));
 sky130_fd_sc_hd__nor2_1 _13108_ (.A(_05856_),
    .B(_05861_),
    .Y(_05888_));
 sky130_fd_sc_hd__nand2_1 _13109_ (.A(\top_inst.grid_inst.data_path_wires[1][1] ),
    .B(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[6] ),
    .Y(_05889_));
 sky130_fd_sc_hd__or2b_1 _13110_ (.A(\top_inst.grid_inst.data_path_wires[1][0] ),
    .B_N(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[7] ),
    .X(_05890_));
 sky130_fd_sc_hd__xnor2_1 _13111_ (.A(_05889_),
    .B(_05890_),
    .Y(_05891_));
 sky130_fd_sc_hd__nand2_1 _13112_ (.A(_05741_),
    .B(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[5] ),
    .Y(_05892_));
 sky130_fd_sc_hd__xnor2_1 _13113_ (.A(_05891_),
    .B(_05892_),
    .Y(_05893_));
 sky130_fd_sc_hd__xor2_1 _13114_ (.A(_05855_),
    .B(_05893_),
    .X(_05894_));
 sky130_fd_sc_hd__a22o_1 _13115_ (.A1(_05744_),
    .A2(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[1][4] ),
    .X(_05895_));
 sky130_fd_sc_hd__nand4_4 _13116_ (.A(\top_inst.grid_inst.data_path_wires[1][4] ),
    .B(_05744_),
    .C(_05765_),
    .D(_05763_),
    .Y(_05896_));
 sky130_fd_sc_hd__a22o_1 _13117_ (.A1(\top_inst.grid_inst.data_path_wires[1][5] ),
    .A2(_05761_),
    .B1(_05895_),
    .B2(_05896_),
    .X(_05897_));
 sky130_fd_sc_hd__nand4_2 _13118_ (.A(_05748_),
    .B(_05761_),
    .C(_05895_),
    .D(_05896_),
    .Y(_05898_));
 sky130_fd_sc_hd__nand2_1 _13119_ (.A(_05897_),
    .B(_05898_),
    .Y(_05899_));
 sky130_fd_sc_hd__xnor2_1 _13120_ (.A(_05894_),
    .B(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__xnor2_1 _13121_ (.A(_05888_),
    .B(_05900_),
    .Y(_05901_));
 sky130_fd_sc_hd__nand2_1 _13122_ (.A(_05858_),
    .B(_05860_),
    .Y(_05902_));
 sky130_fd_sc_hd__a22o_1 _13123_ (.A1(\top_inst.grid_inst.data_path_wires[1][6] ),
    .A2(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[1][7] ),
    .X(_05903_));
 sky130_fd_sc_hd__and3_1 _13124_ (.A(\top_inst.grid_inst.data_path_wires[1][7] ),
    .B(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[1] ),
    .C(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[0] ),
    .X(_05904_));
 sky130_fd_sc_hd__nand2_1 _13125_ (.A(_05750_),
    .B(_05904_),
    .Y(_05905_));
 sky130_fd_sc_hd__and3_1 _13126_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[7] ),
    .B(_05903_),
    .C(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__a21oi_1 _13127_ (.A1(_05903_),
    .A2(_05905_),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[7] ),
    .Y(_05907_));
 sky130_fd_sc_hd__or2_1 _13128_ (.A(_05906_),
    .B(_05907_),
    .X(_05908_));
 sky130_fd_sc_hd__xnor2_1 _13129_ (.A(_05902_),
    .B(_05908_),
    .Y(_05909_));
 sky130_fd_sc_hd__xnor2_1 _13130_ (.A(_05865_),
    .B(_05909_),
    .Y(_05910_));
 sky130_fd_sc_hd__xor2_1 _13131_ (.A(_05901_),
    .B(_05910_),
    .X(_05911_));
 sky130_fd_sc_hd__or2_1 _13132_ (.A(_05853_),
    .B(_05862_),
    .X(_05912_));
 sky130_fd_sc_hd__o21ai_1 _13133_ (.A1(_05863_),
    .A2(_05871_),
    .B1(_05912_),
    .Y(_05913_));
 sky130_fd_sc_hd__xnor2_1 _13134_ (.A(_05911_),
    .B(_05913_),
    .Y(_05914_));
 sky130_fd_sc_hd__a21o_1 _13135_ (.A1(_05832_),
    .A2(_05870_),
    .B1(_05868_),
    .X(_05915_));
 sky130_fd_sc_hd__xnor2_1 _13136_ (.A(_05914_),
    .B(_05915_),
    .Y(_05916_));
 sky130_fd_sc_hd__inv_2 _13137_ (.A(_05872_),
    .Y(_05917_));
 sky130_fd_sc_hd__a21oi_1 _13138_ (.A1(_05852_),
    .A2(_05917_),
    .B1(_05874_),
    .Y(_05918_));
 sky130_fd_sc_hd__xnor2_1 _13139_ (.A(_05916_),
    .B(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__or3_1 _13140_ (.A(net169),
    .B(_05881_),
    .C(_05919_),
    .X(_05920_));
 sky130_fd_sc_hd__o21ai_2 _13141_ (.A1(net169),
    .A2(_05881_),
    .B1(_05919_),
    .Y(_05921_));
 sky130_fd_sc_hd__and2_1 _13142_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[7] ),
    .B(_05326_),
    .X(_05922_));
 sky130_fd_sc_hd__a31o_1 _13143_ (.A1(_05887_),
    .A2(_05920_),
    .A3(_05921_),
    .B1(_05922_),
    .X(_05923_));
 sky130_fd_sc_hd__and2_1 _13144_ (.A(_05886_),
    .B(_05923_),
    .X(_05924_));
 sky130_fd_sc_hd__clkbuf_1 _13145_ (.A(_05924_),
    .X(_00342_));
 sky130_fd_sc_hd__or2b_1 _13146_ (.A(_05918_),
    .B_N(_05916_),
    .X(_05925_));
 sky130_fd_sc_hd__and2b_1 _13147_ (.A_N(\top_inst.grid_inst.data_path_wires[1][1] ),
    .B(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[7] ),
    .X(_05926_));
 sky130_fd_sc_hd__a21oi_1 _13148_ (.A1(_05741_),
    .A2(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[6] ),
    .B1(_05926_),
    .Y(_05927_));
 sky130_fd_sc_hd__and3_1 _13149_ (.A(\top_inst.grid_inst.data_path_wires[1][2] ),
    .B(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[6] ),
    .C(_05926_),
    .X(_05928_));
 sky130_fd_sc_hd__nor2_1 _13150_ (.A(_05927_),
    .B(_05928_),
    .Y(_05929_));
 sky130_fd_sc_hd__nand2_1 _13151_ (.A(_05744_),
    .B(_05768_),
    .Y(_05930_));
 sky130_fd_sc_hd__xnor2_1 _13152_ (.A(_05929_),
    .B(_05930_),
    .Y(_05931_));
 sky130_fd_sc_hd__nor2_1 _13153_ (.A(_05891_),
    .B(_05892_),
    .Y(_05932_));
 sky130_fd_sc_hd__o21ba_1 _13154_ (.A1(_05889_),
    .A2(_05890_),
    .B1_N(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__xnor2_1 _13155_ (.A(_05931_),
    .B(_05933_),
    .Y(_05934_));
 sky130_fd_sc_hd__a22o_1 _13156_ (.A1(\top_inst.grid_inst.data_path_wires[1][4] ),
    .A2(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[1][5] ),
    .X(_05935_));
 sky130_fd_sc_hd__nand4_1 _13157_ (.A(\top_inst.grid_inst.data_path_wires[1][5] ),
    .B(_05746_),
    .C(_05765_),
    .D(_05763_),
    .Y(_05936_));
 sky130_fd_sc_hd__a22oi_1 _13158_ (.A1(_05750_),
    .A2(_05761_),
    .B1(_05935_),
    .B2(_05936_),
    .Y(_05937_));
 sky130_fd_sc_hd__and4_1 _13159_ (.A(_05750_),
    .B(_05761_),
    .C(_05935_),
    .D(_05936_),
    .X(_05938_));
 sky130_fd_sc_hd__or2_1 _13160_ (.A(_05937_),
    .B(_05938_),
    .X(_05939_));
 sky130_fd_sc_hd__xnor2_1 _13161_ (.A(_05934_),
    .B(_05939_),
    .Y(_05940_));
 sky130_fd_sc_hd__and3_1 _13162_ (.A(_05894_),
    .B(_05897_),
    .C(_05898_),
    .X(_05941_));
 sky130_fd_sc_hd__o21ba_1 _13163_ (.A1(_05855_),
    .A2(_05893_),
    .B1_N(_05941_),
    .X(_05942_));
 sky130_fd_sc_hd__xnor2_1 _13164_ (.A(_05940_),
    .B(_05942_),
    .Y(_05943_));
 sky130_fd_sc_hd__and2_1 _13165_ (.A(_05751_),
    .B(_05904_),
    .X(_05944_));
 sky130_fd_sc_hd__o21ai_4 _13166_ (.A1(_05759_),
    .A2(_05757_),
    .B1(\top_inst.grid_inst.data_path_wires[1][7] ),
    .Y(_05945_));
 sky130_fd_sc_hd__or2_1 _13167_ (.A(_05904_),
    .B(_05945_),
    .X(_05946_));
 sky130_fd_sc_hd__a21o_1 _13168_ (.A1(_05896_),
    .A2(_05898_),
    .B1(_05946_),
    .X(_05947_));
 sky130_fd_sc_hd__nand3_1 _13169_ (.A(_05896_),
    .B(_05898_),
    .C(_05946_),
    .Y(_05948_));
 sky130_fd_sc_hd__o211a_1 _13170_ (.A1(_05944_),
    .A2(_05906_),
    .B1(_05947_),
    .C1(_05948_),
    .X(_05949_));
 sky130_fd_sc_hd__nor2_1 _13171_ (.A(_05944_),
    .B(_05906_),
    .Y(_05950_));
 sky130_fd_sc_hd__a21boi_1 _13172_ (.A1(_05947_),
    .A2(_05948_),
    .B1_N(_05950_),
    .Y(_05951_));
 sky130_fd_sc_hd__nor2_1 _13173_ (.A(_05949_),
    .B(_05951_),
    .Y(_05952_));
 sky130_fd_sc_hd__xnor2_1 _13174_ (.A(_05943_),
    .B(_05952_),
    .Y(_05953_));
 sky130_fd_sc_hd__nand2_1 _13175_ (.A(_05888_),
    .B(_05900_),
    .Y(_05954_));
 sky130_fd_sc_hd__o21a_1 _13176_ (.A1(_05901_),
    .A2(_05910_),
    .B1(_05954_),
    .X(_05955_));
 sky130_fd_sc_hd__xnor2_1 _13177_ (.A(_05953_),
    .B(_05955_),
    .Y(_05956_));
 sky130_fd_sc_hd__or2b_1 _13178_ (.A(_05908_),
    .B_N(_05902_),
    .X(_05957_));
 sky130_fd_sc_hd__a21boi_1 _13179_ (.A1(_05865_),
    .A2(_05909_),
    .B1_N(_05957_),
    .Y(_05958_));
 sky130_fd_sc_hd__xnor2_1 _13180_ (.A(_05956_),
    .B(_05958_),
    .Y(_05959_));
 sky130_fd_sc_hd__or2b_1 _13181_ (.A(_05914_),
    .B_N(_05915_),
    .X(_05960_));
 sky130_fd_sc_hd__a21boi_1 _13182_ (.A1(_05911_),
    .A2(_05913_),
    .B1_N(_05960_),
    .Y(_05961_));
 sky130_fd_sc_hd__xnor2_1 _13183_ (.A(_05959_),
    .B(_05961_),
    .Y(_05962_));
 sky130_fd_sc_hd__a21o_1 _13184_ (.A1(_05925_),
    .A2(_05921_),
    .B1(_05962_),
    .X(_05963_));
 sky130_fd_sc_hd__a31oi_1 _13185_ (.A1(_05925_),
    .A2(_05921_),
    .A3(_05962_),
    .B1(_05405_),
    .Y(_05964_));
 sky130_fd_sc_hd__a22o_1 _13186_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[8] ),
    .A2(_05354_),
    .B1(_05963_),
    .B2(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__and2_1 _13187_ (.A(_05886_),
    .B(_05965_),
    .X(_05966_));
 sky130_fd_sc_hd__clkbuf_1 _13188_ (.A(_05966_),
    .X(_00343_));
 sky130_fd_sc_hd__nor2_1 _13189_ (.A(_05959_),
    .B(_05961_),
    .Y(_05967_));
 sky130_fd_sc_hd__inv_2 _13190_ (.A(_05967_),
    .Y(_05968_));
 sky130_fd_sc_hd__and2b_1 _13191_ (.A_N(\top_inst.grid_inst.data_path_wires[1][2] ),
    .B(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[7] ),
    .X(_05969_));
 sky130_fd_sc_hd__a21oi_1 _13192_ (.A1(_05744_),
    .A2(_05770_),
    .B1(_05969_),
    .Y(_05970_));
 sky130_fd_sc_hd__and3_1 _13193_ (.A(_05744_),
    .B(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[6] ),
    .C(_05969_),
    .X(_05971_));
 sky130_fd_sc_hd__nor2_1 _13194_ (.A(_05970_),
    .B(_05971_),
    .Y(_05972_));
 sky130_fd_sc_hd__nand2_1 _13195_ (.A(_05746_),
    .B(_05768_),
    .Y(_05973_));
 sky130_fd_sc_hd__xnor2_1 _13196_ (.A(_05972_),
    .B(_05973_),
    .Y(_05974_));
 sky130_fd_sc_hd__o21ba_1 _13197_ (.A1(_05927_),
    .A2(_05930_),
    .B1_N(_05928_),
    .X(_05975_));
 sky130_fd_sc_hd__xor2_1 _13198_ (.A(_05974_),
    .B(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__a22oi_2 _13199_ (.A1(_05748_),
    .A2(_05765_),
    .B1(_05763_),
    .B2(_05750_),
    .Y(_05977_));
 sky130_fd_sc_hd__and4_1 _13200_ (.A(_05750_),
    .B(\top_inst.grid_inst.data_path_wires[1][5] ),
    .C(_05765_),
    .D(_05763_),
    .X(_05978_));
 sky130_fd_sc_hd__nor2_1 _13201_ (.A(_05977_),
    .B(_05978_),
    .Y(_05979_));
 sky130_fd_sc_hd__nand2_2 _13202_ (.A(_05753_),
    .B(_05761_),
    .Y(_05980_));
 sky130_fd_sc_hd__xor2_1 _13203_ (.A(_05979_),
    .B(_05980_),
    .X(_05981_));
 sky130_fd_sc_hd__xor2_1 _13204_ (.A(_05976_),
    .B(_05981_),
    .X(_05982_));
 sky130_fd_sc_hd__inv_2 _13205_ (.A(_05933_),
    .Y(_05983_));
 sky130_fd_sc_hd__or3b_1 _13206_ (.A(_05937_),
    .B(_05938_),
    .C_N(_05934_),
    .X(_05984_));
 sky130_fd_sc_hd__a21boi_1 _13207_ (.A1(_05931_),
    .A2(_05983_),
    .B1_N(_05984_),
    .Y(_05985_));
 sky130_fd_sc_hd__xnor2_1 _13208_ (.A(_05982_),
    .B(_05985_),
    .Y(_05986_));
 sky130_fd_sc_hd__and4_1 _13209_ (.A(_05748_),
    .B(_05746_),
    .C(_05765_),
    .D(_05763_),
    .X(_05987_));
 sky130_fd_sc_hd__nor2_1 _13210_ (.A(_05987_),
    .B(_05938_),
    .Y(_05988_));
 sky130_fd_sc_hd__nor2_1 _13211_ (.A(_05945_),
    .B(_05988_),
    .Y(_05989_));
 sky130_fd_sc_hd__and2_1 _13212_ (.A(_05945_),
    .B(_05988_),
    .X(_05990_));
 sky130_fd_sc_hd__nor2_1 _13213_ (.A(_05989_),
    .B(_05990_),
    .Y(_05991_));
 sky130_fd_sc_hd__xnor2_1 _13214_ (.A(_05986_),
    .B(_05991_),
    .Y(_05992_));
 sky130_fd_sc_hd__and2b_1 _13215_ (.A_N(_05942_),
    .B(_05940_),
    .X(_05993_));
 sky130_fd_sc_hd__a21oi_1 _13216_ (.A1(_05943_),
    .A2(_05952_),
    .B1(_05993_),
    .Y(_05994_));
 sky130_fd_sc_hd__xnor2_1 _13217_ (.A(_05992_),
    .B(_05994_),
    .Y(_05995_));
 sky130_fd_sc_hd__and3_1 _13218_ (.A(_05896_),
    .B(_05898_),
    .C(_05946_),
    .X(_05996_));
 sky130_fd_sc_hd__o21a_1 _13219_ (.A1(_05950_),
    .A2(_05996_),
    .B1(_05947_),
    .X(_05997_));
 sky130_fd_sc_hd__xnor2_1 _13220_ (.A(_05995_),
    .B(_05997_),
    .Y(_05998_));
 sky130_fd_sc_hd__or2_1 _13221_ (.A(_05953_),
    .B(_05955_),
    .X(_05999_));
 sky130_fd_sc_hd__o21a_1 _13222_ (.A1(_05956_),
    .A2(_05958_),
    .B1(_05999_),
    .X(_06000_));
 sky130_fd_sc_hd__xnor2_1 _13223_ (.A(_05998_),
    .B(_06000_),
    .Y(_06001_));
 sky130_fd_sc_hd__a21o_1 _13224_ (.A1(_05968_),
    .A2(_05963_),
    .B1(_06001_),
    .X(_06002_));
 sky130_fd_sc_hd__nand3_1 _13225_ (.A(_05968_),
    .B(_05963_),
    .C(_06001_),
    .Y(_06003_));
 sky130_fd_sc_hd__a21o_1 _13226_ (.A1(_06002_),
    .A2(_06003_),
    .B1(_05328_),
    .X(_06004_));
 sky130_fd_sc_hd__o211a_1 _13227_ (.A1(net1024),
    .A2(_05788_),
    .B1(_06004_),
    .C1(_05767_),
    .X(_00344_));
 sky130_fd_sc_hd__or2_1 _13228_ (.A(_05998_),
    .B(_06000_),
    .X(_06005_));
 sky130_fd_sc_hd__or2b_1 _13229_ (.A(_05975_),
    .B_N(_05974_),
    .X(_06006_));
 sky130_fd_sc_hd__o21a_1 _13230_ (.A1(_05976_),
    .A2(_05981_),
    .B1(_06006_),
    .X(_06007_));
 sky130_fd_sc_hd__and2b_1 _13231_ (.A_N(\top_inst.grid_inst.data_path_wires[1][3] ),
    .B(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[7] ),
    .X(_06008_));
 sky130_fd_sc_hd__a21oi_1 _13232_ (.A1(_05746_),
    .A2(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[6] ),
    .B1(_06008_),
    .Y(_06009_));
 sky130_fd_sc_hd__and3_1 _13233_ (.A(\top_inst.grid_inst.data_path_wires[1][4] ),
    .B(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[6] ),
    .C(_06008_),
    .X(_06010_));
 sky130_fd_sc_hd__nor2_1 _13234_ (.A(_06009_),
    .B(_06010_),
    .Y(_06011_));
 sky130_fd_sc_hd__nand2_1 _13235_ (.A(\top_inst.grid_inst.data_path_wires[1][5] ),
    .B(_05768_),
    .Y(_06012_));
 sky130_fd_sc_hd__xnor2_1 _13236_ (.A(_06011_),
    .B(_06012_),
    .Y(_06013_));
 sky130_fd_sc_hd__o21ba_1 _13237_ (.A1(_05970_),
    .A2(_05973_),
    .B1_N(_05971_),
    .X(_06014_));
 sky130_fd_sc_hd__xor2_1 _13238_ (.A(_06013_),
    .B(_06014_),
    .X(_06015_));
 sky130_fd_sc_hd__and3_2 _13239_ (.A(\top_inst.grid_inst.data_path_wires[1][7] ),
    .B(_05765_),
    .C(_05763_),
    .X(_06016_));
 sky130_fd_sc_hd__a22oi_1 _13240_ (.A1(_05750_),
    .A2(_05765_),
    .B1(_05763_),
    .B2(\top_inst.grid_inst.data_path_wires[1][7] ),
    .Y(_06017_));
 sky130_fd_sc_hd__a21oi_1 _13241_ (.A1(_05751_),
    .A2(_06016_),
    .B1(_06017_),
    .Y(_06018_));
 sky130_fd_sc_hd__xnor2_1 _13242_ (.A(_05980_),
    .B(_06018_),
    .Y(_06019_));
 sky130_fd_sc_hd__xnor2_1 _13243_ (.A(_06015_),
    .B(_06019_),
    .Y(_06020_));
 sky130_fd_sc_hd__and2b_1 _13244_ (.A_N(_06007_),
    .B(_06020_),
    .X(_06021_));
 sky130_fd_sc_hd__and2b_1 _13245_ (.A_N(_06020_),
    .B(_06007_),
    .X(_06022_));
 sky130_fd_sc_hd__nor2_1 _13246_ (.A(_06021_),
    .B(_06022_),
    .Y(_06023_));
 sky130_fd_sc_hd__o21ba_1 _13247_ (.A1(_05977_),
    .A2(_05980_),
    .B1_N(_05978_),
    .X(_06024_));
 sky130_fd_sc_hd__nor2_1 _13248_ (.A(_05945_),
    .B(_06024_),
    .Y(_06025_));
 sky130_fd_sc_hd__and2_1 _13249_ (.A(_05945_),
    .B(_06024_),
    .X(_06026_));
 sky130_fd_sc_hd__nor2_1 _13250_ (.A(_06025_),
    .B(_06026_),
    .Y(_06027_));
 sky130_fd_sc_hd__xnor2_1 _13251_ (.A(_06023_),
    .B(_06027_),
    .Y(_06028_));
 sky130_fd_sc_hd__and2b_1 _13252_ (.A_N(_05985_),
    .B(_05982_),
    .X(_06029_));
 sky130_fd_sc_hd__a21oi_1 _13253_ (.A1(_05986_),
    .A2(_05991_),
    .B1(_06029_),
    .Y(_06030_));
 sky130_fd_sc_hd__xor2_1 _13254_ (.A(_06028_),
    .B(_06030_),
    .X(_06031_));
 sky130_fd_sc_hd__xnor2_1 _13255_ (.A(_05989_),
    .B(_06031_),
    .Y(_06032_));
 sky130_fd_sc_hd__or2_1 _13256_ (.A(_05992_),
    .B(_05994_),
    .X(_06033_));
 sky130_fd_sc_hd__o21a_1 _13257_ (.A1(_05995_),
    .A2(_05997_),
    .B1(_06033_),
    .X(_06034_));
 sky130_fd_sc_hd__nor2_1 _13258_ (.A(_06032_),
    .B(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__and2_1 _13259_ (.A(_06032_),
    .B(_06034_),
    .X(_06036_));
 sky130_fd_sc_hd__or2_1 _13260_ (.A(_06035_),
    .B(_06036_),
    .X(_06037_));
 sky130_fd_sc_hd__a21o_1 _13261_ (.A1(_06005_),
    .A2(_06002_),
    .B1(_06037_),
    .X(_06038_));
 sky130_fd_sc_hd__a31oi_1 _13262_ (.A1(_06005_),
    .A2(_06002_),
    .A3(_06037_),
    .B1(_05405_),
    .Y(_06039_));
 sky130_fd_sc_hd__a22o_1 _13263_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[10] ),
    .A2(_05354_),
    .B1(_06038_),
    .B2(_06039_),
    .X(_06040_));
 sky130_fd_sc_hd__and2_1 _13264_ (.A(_05886_),
    .B(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__clkbuf_1 _13265_ (.A(_06041_),
    .X(_00345_));
 sky130_fd_sc_hd__inv_2 _13266_ (.A(_06035_),
    .Y(_06042_));
 sky130_fd_sc_hd__and2b_1 _13267_ (.A_N(\top_inst.grid_inst.data_path_wires[1][4] ),
    .B(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[7] ),
    .X(_06043_));
 sky130_fd_sc_hd__a21oi_1 _13268_ (.A1(_05748_),
    .A2(_05770_),
    .B1(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__and3_1 _13269_ (.A(_05748_),
    .B(_05770_),
    .C(_06043_),
    .X(_06045_));
 sky130_fd_sc_hd__nor2_1 _13270_ (.A(_06044_),
    .B(_06045_),
    .Y(_06046_));
 sky130_fd_sc_hd__nand2_1 _13271_ (.A(_05751_),
    .B(_05768_),
    .Y(_06047_));
 sky130_fd_sc_hd__xnor2_1 _13272_ (.A(_06046_),
    .B(_06047_),
    .Y(_06048_));
 sky130_fd_sc_hd__o21ba_1 _13273_ (.A1(_06009_),
    .A2(_06012_),
    .B1_N(_06010_),
    .X(_06049_));
 sky130_fd_sc_hd__xnor2_1 _13274_ (.A(_06048_),
    .B(_06049_),
    .Y(_06050_));
 sky130_fd_sc_hd__o21ai_1 _13275_ (.A1(_05765_),
    .A2(_05763_),
    .B1(_05753_),
    .Y(_06051_));
 sky130_fd_sc_hd__nor3_1 _13276_ (.A(_05980_),
    .B(_06016_),
    .C(_06051_),
    .Y(_06052_));
 sky130_fd_sc_hd__o21a_1 _13277_ (.A1(_06016_),
    .A2(_06051_),
    .B1(_05980_),
    .X(_06053_));
 sky130_fd_sc_hd__nor2_2 _13278_ (.A(_06052_),
    .B(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__or2_1 _13279_ (.A(_06050_),
    .B(_06054_),
    .X(_06055_));
 sky130_fd_sc_hd__nand2_1 _13280_ (.A(_06050_),
    .B(_06054_),
    .Y(_06056_));
 sky130_fd_sc_hd__nand2_1 _13281_ (.A(_06055_),
    .B(_06056_),
    .Y(_06057_));
 sky130_fd_sc_hd__or2b_1 _13282_ (.A(_06013_),
    .B_N(_06014_),
    .X(_06058_));
 sky130_fd_sc_hd__and2b_1 _13283_ (.A_N(_06014_),
    .B(_06013_),
    .X(_06059_));
 sky130_fd_sc_hd__a21oi_1 _13284_ (.A1(_06058_),
    .A2(_06019_),
    .B1(_06059_),
    .Y(_06060_));
 sky130_fd_sc_hd__nor2_1 _13285_ (.A(_06057_),
    .B(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__and2_1 _13286_ (.A(_06057_),
    .B(_06060_),
    .X(_06062_));
 sky130_fd_sc_hd__nor2_1 _13287_ (.A(_06061_),
    .B(_06062_),
    .Y(_06063_));
 sky130_fd_sc_hd__o2bb2a_1 _13288_ (.A1_N(_05751_),
    .A2_N(_06016_),
    .B1(_06017_),
    .B2(_05980_),
    .X(_06064_));
 sky130_fd_sc_hd__nor2_1 _13289_ (.A(_05945_),
    .B(_06064_),
    .Y(_06065_));
 sky130_fd_sc_hd__and2_1 _13290_ (.A(_05945_),
    .B(_06064_),
    .X(_06066_));
 sky130_fd_sc_hd__nor2_1 _13291_ (.A(_06065_),
    .B(_06066_),
    .Y(_06067_));
 sky130_fd_sc_hd__xnor2_1 _13292_ (.A(_06063_),
    .B(_06067_),
    .Y(_06068_));
 sky130_fd_sc_hd__a21oi_1 _13293_ (.A1(_06023_),
    .A2(_06027_),
    .B1(_06021_),
    .Y(_06069_));
 sky130_fd_sc_hd__nor2_1 _13294_ (.A(_06068_),
    .B(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__and2_1 _13295_ (.A(_06068_),
    .B(_06069_),
    .X(_06071_));
 sky130_fd_sc_hd__nor2_1 _13296_ (.A(_06070_),
    .B(_06071_),
    .Y(_06072_));
 sky130_fd_sc_hd__xnor2_1 _13297_ (.A(_06025_),
    .B(_06072_),
    .Y(_06073_));
 sky130_fd_sc_hd__nor2_1 _13298_ (.A(_06028_),
    .B(_06030_),
    .Y(_06074_));
 sky130_fd_sc_hd__a21oi_1 _13299_ (.A1(_05989_),
    .A2(_06031_),
    .B1(_06074_),
    .Y(_06075_));
 sky130_fd_sc_hd__xnor2_1 _13300_ (.A(_06073_),
    .B(_06075_),
    .Y(_06076_));
 sky130_fd_sc_hd__a21o_1 _13301_ (.A1(_06042_),
    .A2(_06038_),
    .B1(_06076_),
    .X(_06077_));
 sky130_fd_sc_hd__nand3_1 _13302_ (.A(_06042_),
    .B(_06038_),
    .C(_06076_),
    .Y(_06078_));
 sky130_fd_sc_hd__a21o_1 _13303_ (.A1(_06077_),
    .A2(_06078_),
    .B1(_05328_),
    .X(_06079_));
 sky130_fd_sc_hd__o211a_1 _13304_ (.A1(net1033),
    .A2(_05788_),
    .B1(_06079_),
    .C1(_05767_),
    .X(_00346_));
 sky130_fd_sc_hd__or2_1 _13305_ (.A(_06073_),
    .B(_06075_),
    .X(_06080_));
 sky130_fd_sc_hd__or2b_1 _13306_ (.A(_06049_),
    .B_N(_06048_),
    .X(_06081_));
 sky130_fd_sc_hd__inv_2 _13307_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[7] ),
    .Y(_06082_));
 sky130_fd_sc_hd__o2bb2a_1 _13308_ (.A1_N(_05751_),
    .A2_N(_05770_),
    .B1(_06082_),
    .B2(_05748_),
    .X(_06083_));
 sky130_fd_sc_hd__and4b_1 _13309_ (.A_N(_05748_),
    .B(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[7] ),
    .C(_05770_),
    .D(_05750_),
    .X(_06084_));
 sky130_fd_sc_hd__nand2_1 _13310_ (.A(_05753_),
    .B(_05768_),
    .Y(_06085_));
 sky130_fd_sc_hd__o21a_1 _13311_ (.A1(_06083_),
    .A2(_06084_),
    .B1(_06085_),
    .X(_06086_));
 sky130_fd_sc_hd__nor2_1 _13312_ (.A(_06083_),
    .B(_06084_),
    .Y(_06087_));
 sky130_fd_sc_hd__and3_1 _13313_ (.A(_05753_),
    .B(_05768_),
    .C(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__nor2_1 _13314_ (.A(_06086_),
    .B(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__o21ba_1 _13315_ (.A1(_06044_),
    .A2(_06047_),
    .B1_N(_06045_),
    .X(_06090_));
 sky130_fd_sc_hd__xnor2_1 _13316_ (.A(_06089_),
    .B(_06090_),
    .Y(_06091_));
 sky130_fd_sc_hd__xnor2_1 _13317_ (.A(_06054_),
    .B(_06091_),
    .Y(_06092_));
 sky130_fd_sc_hd__a21o_1 _13318_ (.A1(_06081_),
    .A2(_06056_),
    .B1(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__nand3_1 _13319_ (.A(_06081_),
    .B(_06056_),
    .C(_06092_),
    .Y(_06094_));
 sky130_fd_sc_hd__nand2_1 _13320_ (.A(_06093_),
    .B(_06094_),
    .Y(_06095_));
 sky130_fd_sc_hd__o21a_1 _13321_ (.A1(_05759_),
    .A2(_05757_),
    .B1(_05753_),
    .X(_06096_));
 sky130_fd_sc_hd__o21ai_2 _13322_ (.A1(_06016_),
    .A2(net182),
    .B1(_06096_),
    .Y(_06097_));
 sky130_fd_sc_hd__or3_2 _13323_ (.A(_06096_),
    .B(_06016_),
    .C(net182),
    .X(_06098_));
 sky130_fd_sc_hd__nand2_2 _13324_ (.A(_06097_),
    .B(_06098_),
    .Y(_06099_));
 sky130_fd_sc_hd__inv_2 _13325_ (.A(_06099_),
    .Y(_06100_));
 sky130_fd_sc_hd__xnor2_1 _13326_ (.A(_06095_),
    .B(_06100_),
    .Y(_06101_));
 sky130_fd_sc_hd__a21oi_1 _13327_ (.A1(_06063_),
    .A2(_06067_),
    .B1(_06061_),
    .Y(_06102_));
 sky130_fd_sc_hd__xnor2_1 _13328_ (.A(_06101_),
    .B(_06102_),
    .Y(_06103_));
 sky130_fd_sc_hd__xnor2_1 _13329_ (.A(_06065_),
    .B(_06103_),
    .Y(_06104_));
 sky130_fd_sc_hd__a21oi_1 _13330_ (.A1(_06025_),
    .A2(_06072_),
    .B1(_06070_),
    .Y(_06105_));
 sky130_fd_sc_hd__or2_1 _13331_ (.A(_06104_),
    .B(_06105_),
    .X(_06106_));
 sky130_fd_sc_hd__nand2_1 _13332_ (.A(_06104_),
    .B(_06105_),
    .Y(_06107_));
 sky130_fd_sc_hd__nand2_1 _13333_ (.A(_06106_),
    .B(_06107_),
    .Y(_06108_));
 sky130_fd_sc_hd__a21o_1 _13334_ (.A1(_06080_),
    .A2(_06077_),
    .B1(_06108_),
    .X(_06109_));
 sky130_fd_sc_hd__a31oi_1 _13335_ (.A1(_06080_),
    .A2(_06077_),
    .A3(_06108_),
    .B1(_05405_),
    .Y(_06110_));
 sky130_fd_sc_hd__a22o_1 _13336_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[12] ),
    .A2(_05354_),
    .B1(_06109_),
    .B2(_06110_),
    .X(_06111_));
 sky130_fd_sc_hd__and2_1 _13337_ (.A(_05886_),
    .B(_06111_),
    .X(_06112_));
 sky130_fd_sc_hd__clkbuf_1 _13338_ (.A(_06112_),
    .X(_00347_));
 sky130_fd_sc_hd__inv_2 _13339_ (.A(_06097_),
    .Y(_06113_));
 sky130_fd_sc_hd__o21a_1 _13340_ (.A1(_06095_),
    .A2(_06099_),
    .B1(_06093_),
    .X(_06114_));
 sky130_fd_sc_hd__nand2_1 _13341_ (.A(\top_inst.grid_inst.data_path_wires[1][7] ),
    .B(_05770_),
    .Y(_06115_));
 sky130_fd_sc_hd__o21a_1 _13342_ (.A1(_05751_),
    .A2(_06082_),
    .B1(_06115_),
    .X(_06116_));
 sky130_fd_sc_hd__nor3_1 _13343_ (.A(_05751_),
    .B(_06082_),
    .C(_06115_),
    .Y(_06117_));
 sky130_fd_sc_hd__nor2_1 _13344_ (.A(_06116_),
    .B(_06117_),
    .Y(_06118_));
 sky130_fd_sc_hd__xnor2_1 _13345_ (.A(_06085_),
    .B(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__o21ai_1 _13346_ (.A1(_06084_),
    .A2(_06088_),
    .B1(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__or3_1 _13347_ (.A(_06084_),
    .B(_06088_),
    .C(_06119_),
    .X(_06121_));
 sky130_fd_sc_hd__and2_1 _13348_ (.A(_06120_),
    .B(_06121_),
    .X(_06122_));
 sky130_fd_sc_hd__nand2_1 _13349_ (.A(_06054_),
    .B(_06122_),
    .Y(_06123_));
 sky130_fd_sc_hd__or2_1 _13350_ (.A(_06054_),
    .B(_06122_),
    .X(_06124_));
 sky130_fd_sc_hd__nand2_1 _13351_ (.A(_06123_),
    .B(_06124_),
    .Y(_06125_));
 sky130_fd_sc_hd__or2b_1 _13352_ (.A(_06090_),
    .B_N(_06089_),
    .X(_06126_));
 sky130_fd_sc_hd__a21bo_1 _13353_ (.A1(_06054_),
    .A2(_06091_),
    .B1_N(_06126_),
    .X(_06127_));
 sky130_fd_sc_hd__xor2_1 _13354_ (.A(_06125_),
    .B(_06127_),
    .X(_06128_));
 sky130_fd_sc_hd__xnor2_1 _13355_ (.A(_06100_),
    .B(_06128_),
    .Y(_06129_));
 sky130_fd_sc_hd__and2b_1 _13356_ (.A_N(_06114_),
    .B(_06129_),
    .X(_06130_));
 sky130_fd_sc_hd__and2b_1 _13357_ (.A_N(_06129_),
    .B(_06114_),
    .X(_06131_));
 sky130_fd_sc_hd__nor2_1 _13358_ (.A(_06130_),
    .B(_06131_),
    .Y(_06132_));
 sky130_fd_sc_hd__xnor2_1 _13359_ (.A(_06113_),
    .B(_06132_),
    .Y(_06133_));
 sky130_fd_sc_hd__and2b_1 _13360_ (.A_N(_06102_),
    .B(_06101_),
    .X(_06134_));
 sky130_fd_sc_hd__a21oi_1 _13361_ (.A1(_06065_),
    .A2(_06103_),
    .B1(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__or2_1 _13362_ (.A(_06133_),
    .B(_06135_),
    .X(_06136_));
 sky130_fd_sc_hd__nand2_1 _13363_ (.A(_06133_),
    .B(_06135_),
    .Y(_06137_));
 sky130_fd_sc_hd__nand2_1 _13364_ (.A(_06136_),
    .B(_06137_),
    .Y(_06138_));
 sky130_fd_sc_hd__and3_1 _13365_ (.A(_06106_),
    .B(_06109_),
    .C(_06138_),
    .X(_06139_));
 sky130_fd_sc_hd__clkbuf_16 _13366_ (.A(_05311_),
    .X(_06140_));
 sky130_fd_sc_hd__a21o_1 _13367_ (.A1(_06106_),
    .A2(_06109_),
    .B1(_06138_),
    .X(_06141_));
 sky130_fd_sc_hd__nand2_1 _13368_ (.A(_06140_),
    .B(_06141_),
    .Y(_06142_));
 sky130_fd_sc_hd__a2bb2o_1 _13369_ (.A1_N(_06139_),
    .A2_N(_06142_),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[13] ),
    .B2(_05327_),
    .X(_06143_));
 sky130_fd_sc_hd__and2_1 _13370_ (.A(_05886_),
    .B(_06143_),
    .X(_06144_));
 sky130_fd_sc_hd__clkbuf_1 _13371_ (.A(_06144_),
    .X(_00348_));
 sky130_fd_sc_hd__or2b_1 _13372_ (.A(_06125_),
    .B_N(_06127_),
    .X(_06145_));
 sky130_fd_sc_hd__o21a_1 _13373_ (.A1(_06099_),
    .A2(_06128_),
    .B1(_06145_),
    .X(_06146_));
 sky130_fd_sc_hd__and3_1 _13374_ (.A(_05753_),
    .B(_05770_),
    .C(_05768_),
    .X(_06147_));
 sky130_fd_sc_hd__o21ba_1 _13375_ (.A1(_06085_),
    .A2(_06116_),
    .B1_N(_06117_),
    .X(_06148_));
 sky130_fd_sc_hd__o211a_1 _13376_ (.A1(_05753_),
    .A2(_06082_),
    .B1(_06085_),
    .C1(_06115_),
    .X(_06149_));
 sky130_fd_sc_hd__o21ba_1 _13377_ (.A1(_06147_),
    .A2(_06148_),
    .B1_N(_06149_),
    .X(_06150_));
 sky130_fd_sc_hd__xnor2_1 _13378_ (.A(_06054_),
    .B(_06150_),
    .Y(_06151_));
 sky130_fd_sc_hd__a21oi_1 _13379_ (.A1(_06120_),
    .A2(_06123_),
    .B1(_06151_),
    .Y(_06152_));
 sky130_fd_sc_hd__and3_1 _13380_ (.A(_06120_),
    .B(_06123_),
    .C(_06151_),
    .X(_06153_));
 sky130_fd_sc_hd__nor2_1 _13381_ (.A(_06152_),
    .B(_06153_),
    .Y(_06154_));
 sky130_fd_sc_hd__xnor2_1 _13382_ (.A(_06099_),
    .B(_06154_),
    .Y(_06155_));
 sky130_fd_sc_hd__and2b_1 _13383_ (.A_N(_06146_),
    .B(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__and2b_1 _13384_ (.A_N(_06155_),
    .B(_06146_),
    .X(_06157_));
 sky130_fd_sc_hd__nor2_1 _13385_ (.A(_06156_),
    .B(_06157_),
    .Y(_06158_));
 sky130_fd_sc_hd__xnor2_1 _13386_ (.A(_06113_),
    .B(_06158_),
    .Y(_06159_));
 sky130_fd_sc_hd__a21oi_1 _13387_ (.A1(_06113_),
    .A2(_06132_),
    .B1(_06130_),
    .Y(_06160_));
 sky130_fd_sc_hd__or2_1 _13388_ (.A(_06159_),
    .B(_06160_),
    .X(_06161_));
 sky130_fd_sc_hd__nand2_1 _13389_ (.A(_06159_),
    .B(_06160_),
    .Y(_06162_));
 sky130_fd_sc_hd__nand2_1 _13390_ (.A(_06161_),
    .B(_06162_),
    .Y(_06163_));
 sky130_fd_sc_hd__a21o_1 _13391_ (.A1(_06136_),
    .A2(_06141_),
    .B1(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__a31oi_1 _13392_ (.A1(_06136_),
    .A2(_06141_),
    .A3(_06163_),
    .B1(_05405_),
    .Y(_06165_));
 sky130_fd_sc_hd__a22o_1 _13393_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[14] ),
    .A2(_05354_),
    .B1(_06164_),
    .B2(_06165_),
    .X(_06166_));
 sky130_fd_sc_hd__and2_1 _13394_ (.A(_05886_),
    .B(_06166_),
    .X(_06167_));
 sky130_fd_sc_hd__clkbuf_1 _13395_ (.A(_06167_),
    .X(_00349_));
 sky130_fd_sc_hd__buf_8 _13396_ (.A(_05312_),
    .X(_06168_));
 sky130_fd_sc_hd__buf_8 _13397_ (.A(_06168_),
    .X(_06169_));
 sky130_fd_sc_hd__and3_1 _13398_ (.A(_06098_),
    .B(_06161_),
    .C(_06164_),
    .X(_06170_));
 sky130_fd_sc_hd__a21oi_1 _13399_ (.A1(_06161_),
    .A2(_06164_),
    .B1(_06098_),
    .Y(_06171_));
 sky130_fd_sc_hd__nor2_1 _13400_ (.A(_06054_),
    .B(_06150_),
    .Y(_06172_));
 sky130_fd_sc_hd__a21oi_1 _13401_ (.A1(_06113_),
    .A2(_06158_),
    .B1(_06156_),
    .Y(_06173_));
 sky130_fd_sc_hd__a21oi_1 _13402_ (.A1(_06100_),
    .A2(_06154_),
    .B1(_06152_),
    .Y(_06174_));
 sky130_fd_sc_hd__xnor2_1 _13403_ (.A(_06173_),
    .B(_06174_),
    .Y(_06175_));
 sky130_fd_sc_hd__xnor2_1 _13404_ (.A(_06172_),
    .B(_06175_),
    .Y(_06176_));
 sky130_fd_sc_hd__o21a_1 _13405_ (.A1(_06170_),
    .A2(_06171_),
    .B1(_06176_),
    .X(_06177_));
 sky130_fd_sc_hd__buf_12 _13406_ (.A(_05335_),
    .X(_06178_));
 sky130_fd_sc_hd__o31ai_1 _13407_ (.A1(_06170_),
    .A2(_06171_),
    .A3(_06176_),
    .B1(_06178_),
    .Y(_06179_));
 sky130_fd_sc_hd__clkbuf_16 _13408_ (.A(_04874_),
    .X(_06180_));
 sky130_fd_sc_hd__o221a_1 _13409_ (.A1(net1035),
    .A2(_06169_),
    .B1(_06177_),
    .B2(_06179_),
    .C1(_06180_),
    .X(_00350_));
 sky130_fd_sc_hd__clkbuf_4 _13410_ (.A(\top_inst.grid_inst.data_path_wires[2][0] ),
    .X(_06181_));
 sky130_fd_sc_hd__or2_1 _13411_ (.A(_06181_),
    .B(_05262_),
    .X(_06182_));
 sky130_fd_sc_hd__buf_2 _13412_ (.A(_05260_),
    .X(_06183_));
 sky130_fd_sc_hd__o211a_1 _13413_ (.A1(_05734_),
    .A2(_05256_),
    .B1(_06182_),
    .C1(_06183_),
    .X(_00351_));
 sky130_fd_sc_hd__clkbuf_4 _13414_ (.A(\top_inst.grid_inst.data_path_wires[2][1] ),
    .X(_06184_));
 sky130_fd_sc_hd__or2_1 _13415_ (.A(_06184_),
    .B(_05262_),
    .X(_06185_));
 sky130_fd_sc_hd__o211a_1 _13416_ (.A1(_05738_),
    .A2(_05256_),
    .B1(_06185_),
    .C1(_06183_),
    .X(_00352_));
 sky130_fd_sc_hd__clkbuf_4 _13417_ (.A(\top_inst.grid_inst.data_path_wires[2][2] ),
    .X(_06186_));
 sky130_fd_sc_hd__or2_1 _13418_ (.A(_06186_),
    .B(_05262_),
    .X(_06187_));
 sky130_fd_sc_hd__o211a_1 _13419_ (.A1(_05741_),
    .A2(_05256_),
    .B1(_06187_),
    .C1(_06183_),
    .X(_00353_));
 sky130_fd_sc_hd__buf_4 _13420_ (.A(\top_inst.grid_inst.data_path_wires[2][3] ),
    .X(_06188_));
 sky130_fd_sc_hd__or2_1 _13421_ (.A(_06188_),
    .B(_05262_),
    .X(_06189_));
 sky130_fd_sc_hd__o211a_1 _13422_ (.A1(_05744_),
    .A2(_05256_),
    .B1(_06189_),
    .C1(_06183_),
    .X(_00354_));
 sky130_fd_sc_hd__clkbuf_4 _13423_ (.A(\top_inst.grid_inst.data_path_wires[2][4] ),
    .X(_06190_));
 sky130_fd_sc_hd__or2_1 _13424_ (.A(_06190_),
    .B(_05262_),
    .X(_06191_));
 sky130_fd_sc_hd__o211a_1 _13425_ (.A1(_05746_),
    .A2(_05256_),
    .B1(_06191_),
    .C1(_06183_),
    .X(_00355_));
 sky130_fd_sc_hd__clkbuf_4 _13426_ (.A(_05177_),
    .X(_06192_));
 sky130_fd_sc_hd__buf_4 _13427_ (.A(\top_inst.grid_inst.data_path_wires[2][5] ),
    .X(_06193_));
 sky130_fd_sc_hd__or2_1 _13428_ (.A(_06193_),
    .B(_05262_),
    .X(_06194_));
 sky130_fd_sc_hd__o211a_1 _13429_ (.A1(_05748_),
    .A2(_06192_),
    .B1(_06194_),
    .C1(_06183_),
    .X(_00356_));
 sky130_fd_sc_hd__buf_2 _13430_ (.A(\top_inst.grid_inst.data_path_wires[2][6] ),
    .X(_06195_));
 sky130_fd_sc_hd__clkbuf_4 _13431_ (.A(_06195_),
    .X(_06196_));
 sky130_fd_sc_hd__or2_1 _13432_ (.A(_06196_),
    .B(_05262_),
    .X(_06197_));
 sky130_fd_sc_hd__o211a_1 _13433_ (.A1(_05751_),
    .A2(_06192_),
    .B1(_06197_),
    .C1(_06183_),
    .X(_00357_));
 sky130_fd_sc_hd__clkbuf_4 _13434_ (.A(\top_inst.grid_inst.data_path_wires[2][7] ),
    .X(_06198_));
 sky130_fd_sc_hd__or2_1 _13435_ (.A(_06198_),
    .B(_05262_),
    .X(_06199_));
 sky130_fd_sc_hd__o211a_1 _13436_ (.A1(_05753_),
    .A2(_06192_),
    .B1(_06199_),
    .C1(_06183_),
    .X(_00358_));
 sky130_fd_sc_hd__clkbuf_4 _13437_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[0] ),
    .X(_06200_));
 sky130_fd_sc_hd__or2_1 _13438_ (.A(_06200_),
    .B(_05773_),
    .X(_06201_));
 sky130_fd_sc_hd__o211a_1 _13439_ (.A1(_06181_),
    .A2(_05756_),
    .B1(_06201_),
    .C1(_06183_),
    .X(_00359_));
 sky130_fd_sc_hd__clkbuf_4 _13440_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[1] ),
    .X(_06202_));
 sky130_fd_sc_hd__or2_1 _13441_ (.A(_06202_),
    .B(_05773_),
    .X(_06203_));
 sky130_fd_sc_hd__o211a_1 _13442_ (.A1(_06184_),
    .A2(_05756_),
    .B1(_06203_),
    .C1(_06183_),
    .X(_00360_));
 sky130_fd_sc_hd__clkbuf_4 _13443_ (.A(_05755_),
    .X(_06204_));
 sky130_fd_sc_hd__clkbuf_4 _13444_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[2] ),
    .X(_06205_));
 sky130_fd_sc_hd__or2_1 _13445_ (.A(_06205_),
    .B(_05773_),
    .X(_06206_));
 sky130_fd_sc_hd__clkbuf_4 _13446_ (.A(_05260_),
    .X(_06207_));
 sky130_fd_sc_hd__o211a_1 _13447_ (.A1(_06186_),
    .A2(_06204_),
    .B1(_06206_),
    .C1(_06207_),
    .X(_00361_));
 sky130_fd_sc_hd__clkbuf_4 _13448_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[3] ),
    .X(_06208_));
 sky130_fd_sc_hd__or2_1 _13449_ (.A(_06208_),
    .B(_05773_),
    .X(_06209_));
 sky130_fd_sc_hd__o211a_1 _13450_ (.A1(_06188_),
    .A2(_06204_),
    .B1(_06209_),
    .C1(_06207_),
    .X(_00362_));
 sky130_fd_sc_hd__clkbuf_4 _13451_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[4] ),
    .X(_06210_));
 sky130_fd_sc_hd__or2_1 _13452_ (.A(_06210_),
    .B(_05773_),
    .X(_06211_));
 sky130_fd_sc_hd__o211a_1 _13453_ (.A1(_06190_),
    .A2(_06204_),
    .B1(_06211_),
    .C1(_06207_),
    .X(_00363_));
 sky130_fd_sc_hd__clkbuf_4 _13454_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[5] ),
    .X(_06212_));
 sky130_fd_sc_hd__or2_1 _13455_ (.A(_06212_),
    .B(_05773_),
    .X(_06213_));
 sky130_fd_sc_hd__o211a_1 _13456_ (.A1(_06193_),
    .A2(_06204_),
    .B1(_06213_),
    .C1(_06207_),
    .X(_00364_));
 sky130_fd_sc_hd__buf_2 _13457_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[6] ),
    .X(_06214_));
 sky130_fd_sc_hd__or2_1 _13458_ (.A(_06214_),
    .B(_05773_),
    .X(_06215_));
 sky130_fd_sc_hd__o211a_1 _13459_ (.A1(_06196_),
    .A2(_06204_),
    .B1(_06215_),
    .C1(_06207_),
    .X(_00365_));
 sky130_fd_sc_hd__or2_1 _13460_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[7] ),
    .B(_05773_),
    .X(_06216_));
 sky130_fd_sc_hd__o211a_1 _13461_ (.A1(_06198_),
    .A2(_06204_),
    .B1(_06216_),
    .C1(_06207_),
    .X(_00366_));
 sky130_fd_sc_hd__nand2_1 _13462_ (.A(_06181_),
    .B(_06200_),
    .Y(_06217_));
 sky130_fd_sc_hd__nand2_1 _13463_ (.A(_05317_),
    .B(_06217_),
    .Y(_06218_));
 sky130_fd_sc_hd__o211a_1 _13464_ (.A1(net1017),
    .A2(_05788_),
    .B1(_06218_),
    .C1(_06207_),
    .X(_00367_));
 sky130_fd_sc_hd__nand2_1 _13465_ (.A(_06184_),
    .B(_06202_),
    .Y(_06219_));
 sky130_fd_sc_hd__a22o_1 _13466_ (.A1(_06181_),
    .A2(_06202_),
    .B1(_06200_),
    .B2(_06184_),
    .X(_06220_));
 sky130_fd_sc_hd__o21ai_1 _13467_ (.A1(_06217_),
    .A2(_06219_),
    .B1(_06220_),
    .Y(_06221_));
 sky130_fd_sc_hd__nand2_1 _13468_ (.A(_05317_),
    .B(_06221_),
    .Y(_06222_));
 sky130_fd_sc_hd__o211a_1 _13469_ (.A1(net1004),
    .A2(_05788_),
    .B1(_06222_),
    .C1(_06207_),
    .X(_00368_));
 sky130_fd_sc_hd__nand2_1 _13470_ (.A(_06186_),
    .B(_06200_),
    .Y(_06223_));
 sky130_fd_sc_hd__and3_1 _13471_ (.A(_06184_),
    .B(_06202_),
    .C(_06217_),
    .X(_06224_));
 sky130_fd_sc_hd__xnor2_1 _13472_ (.A(_06223_),
    .B(_06224_),
    .Y(_06225_));
 sky130_fd_sc_hd__a21oi_1 _13473_ (.A1(_06181_),
    .A2(_06205_),
    .B1(_06225_),
    .Y(_06226_));
 sky130_fd_sc_hd__and3_1 _13474_ (.A(_06181_),
    .B(_06205_),
    .C(_06225_),
    .X(_06227_));
 sky130_fd_sc_hd__o21ai_1 _13475_ (.A1(_06226_),
    .A2(_06227_),
    .B1(_05336_),
    .Y(_06228_));
 sky130_fd_sc_hd__o211a_1 _13476_ (.A1(net1056),
    .A2(_05788_),
    .B1(_06228_),
    .C1(_06207_),
    .X(_00369_));
 sky130_fd_sc_hd__a22oi_1 _13477_ (.A1(_06181_),
    .A2(_06208_),
    .B1(_06205_),
    .B2(_06184_),
    .Y(_06229_));
 sky130_fd_sc_hd__and4_1 _13478_ (.A(\top_inst.grid_inst.data_path_wires[2][1] ),
    .B(\top_inst.grid_inst.data_path_wires[2][0] ),
    .C(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[3] ),
    .D(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[2] ),
    .X(_06230_));
 sky130_fd_sc_hd__or2_1 _13479_ (.A(_06229_),
    .B(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__and4_1 _13480_ (.A(\top_inst.grid_inst.data_path_wires[2][3] ),
    .B(\top_inst.grid_inst.data_path_wires[2][2] ),
    .C(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[0] ),
    .X(_06232_));
 sky130_fd_sc_hd__o21a_1 _13481_ (.A1(_06219_),
    .A2(_06223_),
    .B1(_06232_),
    .X(_06233_));
 sky130_fd_sc_hd__a22o_1 _13482_ (.A1(_06186_),
    .A2(_06202_),
    .B1(_06200_),
    .B2(_06188_),
    .X(_06234_));
 sky130_fd_sc_hd__or3_2 _13483_ (.A(_06219_),
    .B(_06223_),
    .C(_06232_),
    .X(_06235_));
 sky130_fd_sc_hd__and3b_1 _13484_ (.A_N(_06233_),
    .B(_06234_),
    .C(_06235_),
    .X(_06236_));
 sky130_fd_sc_hd__xnor2_1 _13485_ (.A(_06231_),
    .B(_06236_),
    .Y(_06237_));
 sky130_fd_sc_hd__nor3_1 _13486_ (.A(_06186_),
    .B(_06217_),
    .C(_06219_),
    .Y(_06238_));
 sky130_fd_sc_hd__nor3_1 _13487_ (.A(_06227_),
    .B(_06237_),
    .C(_06238_),
    .Y(_06239_));
 sky130_fd_sc_hd__o21a_1 _13488_ (.A1(_06227_),
    .A2(_06238_),
    .B1(_06237_),
    .X(_06240_));
 sky130_fd_sc_hd__o21ai_1 _13489_ (.A1(_06239_),
    .A2(_06240_),
    .B1(_05336_),
    .Y(_06241_));
 sky130_fd_sc_hd__o211a_1 _13490_ (.A1(net1031),
    .A2(_05788_),
    .B1(_06241_),
    .C1(_06207_),
    .X(_00370_));
 sky130_fd_sc_hd__clkbuf_8 _13491_ (.A(_05353_),
    .X(_06242_));
 sky130_fd_sc_hd__and2b_1 _13492_ (.A_N(_06231_),
    .B(_06236_),
    .X(_06243_));
 sky130_fd_sc_hd__inv_2 _13493_ (.A(_06232_),
    .Y(_06244_));
 sky130_fd_sc_hd__nand4_1 _13494_ (.A(\top_inst.grid_inst.data_path_wires[2][4] ),
    .B(\top_inst.grid_inst.data_path_wires[2][3] ),
    .C(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[0] ),
    .Y(_06245_));
 sky130_fd_sc_hd__a22o_1 _13495_ (.A1(\top_inst.grid_inst.data_path_wires[2][3] ),
    .A2(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[2][4] ),
    .X(_06246_));
 sky130_fd_sc_hd__and3_1 _13496_ (.A(_06230_),
    .B(_06245_),
    .C(_06246_),
    .X(_06247_));
 sky130_fd_sc_hd__a21oi_1 _13497_ (.A1(_06245_),
    .A2(_06246_),
    .B1(_06230_),
    .Y(_06248_));
 sky130_fd_sc_hd__nor2_1 _13498_ (.A(_06247_),
    .B(_06248_),
    .Y(_06249_));
 sky130_fd_sc_hd__xnor2_1 _13499_ (.A(_06244_),
    .B(_06249_),
    .Y(_06250_));
 sky130_fd_sc_hd__nand2_1 _13500_ (.A(_06186_),
    .B(_06205_),
    .Y(_06251_));
 sky130_fd_sc_hd__and3_1 _13501_ (.A(\top_inst.grid_inst.data_path_wires[2][1] ),
    .B(\top_inst.grid_inst.data_path_wires[2][0] ),
    .C(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[3] ),
    .X(_06252_));
 sky130_fd_sc_hd__a22o_1 _13502_ (.A1(\top_inst.grid_inst.data_path_wires[2][0] ),
    .A2(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[2][1] ),
    .X(_06253_));
 sky130_fd_sc_hd__a21bo_1 _13503_ (.A1(_06210_),
    .A2(_06252_),
    .B1_N(_06253_),
    .X(_06254_));
 sky130_fd_sc_hd__xor2_1 _13504_ (.A(_06251_),
    .B(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__xor2_1 _13505_ (.A(_06250_),
    .B(_06255_),
    .X(_06256_));
 sky130_fd_sc_hd__xnor2_1 _13506_ (.A(_06243_),
    .B(_06256_),
    .Y(_06257_));
 sky130_fd_sc_hd__xor2_1 _13507_ (.A(_06235_),
    .B(_06257_),
    .X(_06258_));
 sky130_fd_sc_hd__nand2_1 _13508_ (.A(_06240_),
    .B(_06258_),
    .Y(_06259_));
 sky130_fd_sc_hd__o21a_1 _13509_ (.A1(_06240_),
    .A2(_06258_),
    .B1(_05315_),
    .X(_06260_));
 sky130_fd_sc_hd__a22o_1 _13510_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[4] ),
    .A2(_06242_),
    .B1(_06259_),
    .B2(_06260_),
    .X(_06261_));
 sky130_fd_sc_hd__and2_1 _13511_ (.A(_05886_),
    .B(_06261_),
    .X(_06262_));
 sky130_fd_sc_hd__clkbuf_1 _13512_ (.A(_06262_),
    .X(_00371_));
 sky130_fd_sc_hd__and2_1 _13513_ (.A(_06250_),
    .B(_06255_),
    .X(_06263_));
 sky130_fd_sc_hd__nand2_1 _13514_ (.A(_06181_),
    .B(_06212_),
    .Y(_06264_));
 sky130_fd_sc_hd__a22o_1 _13515_ (.A1(\top_inst.grid_inst.data_path_wires[2][1] ),
    .A2(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[2][2] ),
    .X(_06265_));
 sky130_fd_sc_hd__nand4_1 _13516_ (.A(\top_inst.grid_inst.data_path_wires[2][2] ),
    .B(_06184_),
    .C(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[3] ),
    .Y(_06266_));
 sky130_fd_sc_hd__nand2_1 _13517_ (.A(_06265_),
    .B(_06266_),
    .Y(_06267_));
 sky130_fd_sc_hd__and2_1 _13518_ (.A(\top_inst.grid_inst.data_path_wires[2][3] ),
    .B(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[2] ),
    .X(_06268_));
 sky130_fd_sc_hd__xor2_2 _13519_ (.A(_06267_),
    .B(_06268_),
    .X(_06269_));
 sky130_fd_sc_hd__xor2_2 _13520_ (.A(_06264_),
    .B(_06269_),
    .X(_06270_));
 sky130_fd_sc_hd__and4_1 _13521_ (.A(_06190_),
    .B(_06188_),
    .C(_06202_),
    .D(_06200_),
    .X(_06271_));
 sky130_fd_sc_hd__a32o_1 _13522_ (.A1(\top_inst.grid_inst.data_path_wires[2][2] ),
    .A2(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[2] ),
    .A3(_06253_),
    .B1(_06252_),
    .B2(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[4] ),
    .X(_06272_));
 sky130_fd_sc_hd__and4_2 _13523_ (.A(\top_inst.grid_inst.data_path_wires[2][5] ),
    .B(\top_inst.grid_inst.data_path_wires[2][4] ),
    .C(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[0] ),
    .X(_06273_));
 sky130_fd_sc_hd__a22oi_1 _13524_ (.A1(\top_inst.grid_inst.data_path_wires[2][4] ),
    .A2(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[2][5] ),
    .Y(_06274_));
 sky130_fd_sc_hd__nor2_1 _13525_ (.A(_06273_),
    .B(_06274_),
    .Y(_06275_));
 sky130_fd_sc_hd__xor2_2 _13526_ (.A(_06272_),
    .B(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__xnor2_2 _13527_ (.A(_06271_),
    .B(_06276_),
    .Y(_06277_));
 sky130_fd_sc_hd__xor2_2 _13528_ (.A(_06270_),
    .B(_06277_),
    .X(_06278_));
 sky130_fd_sc_hd__xnor2_1 _13529_ (.A(_06263_),
    .B(_06278_),
    .Y(_06279_));
 sky130_fd_sc_hd__o21ba_1 _13530_ (.A1(_06244_),
    .A2(_06248_),
    .B1_N(_06247_),
    .X(_06280_));
 sky130_fd_sc_hd__xor2_1 _13531_ (.A(_06279_),
    .B(_06280_),
    .X(_06281_));
 sky130_fd_sc_hd__nand2_1 _13532_ (.A(_06243_),
    .B(_06256_),
    .Y(_06282_));
 sky130_fd_sc_hd__o21a_1 _13533_ (.A1(_06235_),
    .A2(_06257_),
    .B1(_06282_),
    .X(_06283_));
 sky130_fd_sc_hd__xnor2_1 _13534_ (.A(_06281_),
    .B(_06283_),
    .Y(_06284_));
 sky130_fd_sc_hd__or2_1 _13535_ (.A(_06259_),
    .B(_06284_),
    .X(_06285_));
 sky130_fd_sc_hd__a21oi_1 _13536_ (.A1(_06259_),
    .A2(_06284_),
    .B1(_05399_),
    .Y(_06286_));
 sky130_fd_sc_hd__a22o_1 _13537_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[5] ),
    .A2(_06242_),
    .B1(_06285_),
    .B2(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__and2_1 _13538_ (.A(_05886_),
    .B(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__clkbuf_1 _13539_ (.A(_06288_),
    .X(_00372_));
 sky130_fd_sc_hd__or2_1 _13540_ (.A(_06281_),
    .B(_06283_),
    .X(_06289_));
 sky130_fd_sc_hd__nand2_1 _13541_ (.A(_06272_),
    .B(_06275_),
    .Y(_06290_));
 sky130_fd_sc_hd__nand2_1 _13542_ (.A(_06271_),
    .B(_06276_),
    .Y(_06291_));
 sky130_fd_sc_hd__inv_2 _13543_ (.A(_06270_),
    .Y(_06292_));
 sky130_fd_sc_hd__nor2_1 _13544_ (.A(_06292_),
    .B(_06277_),
    .Y(_06293_));
 sky130_fd_sc_hd__or2_1 _13545_ (.A(_06264_),
    .B(_06269_),
    .X(_06294_));
 sky130_fd_sc_hd__a22o_1 _13546_ (.A1(_06181_),
    .A2(_06214_),
    .B1(_06212_),
    .B2(_06184_),
    .X(_06295_));
 sky130_fd_sc_hd__nand4_2 _13547_ (.A(_06184_),
    .B(\top_inst.grid_inst.data_path_wires[2][0] ),
    .C(_06214_),
    .D(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[5] ),
    .Y(_06296_));
 sky130_fd_sc_hd__nand2_1 _13548_ (.A(_06295_),
    .B(_06296_),
    .Y(_06297_));
 sky130_fd_sc_hd__a22o_1 _13549_ (.A1(\top_inst.grid_inst.data_path_wires[2][2] ),
    .A2(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[2][3] ),
    .X(_06298_));
 sky130_fd_sc_hd__nand4_2 _13550_ (.A(\top_inst.grid_inst.data_path_wires[2][3] ),
    .B(_06186_),
    .C(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[3] ),
    .Y(_06299_));
 sky130_fd_sc_hd__a22o_1 _13551_ (.A1(_06190_),
    .A2(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[2] ),
    .B1(_06298_),
    .B2(_06299_),
    .X(_06300_));
 sky130_fd_sc_hd__nand4_1 _13552_ (.A(_06190_),
    .B(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[2] ),
    .C(_06298_),
    .D(_06299_),
    .Y(_06301_));
 sky130_fd_sc_hd__nand2_1 _13553_ (.A(_06300_),
    .B(_06301_),
    .Y(_06302_));
 sky130_fd_sc_hd__xnor2_2 _13554_ (.A(_06297_),
    .B(_06302_),
    .Y(_06303_));
 sky130_fd_sc_hd__xnor2_2 _13555_ (.A(_06294_),
    .B(_06303_),
    .Y(_06304_));
 sky130_fd_sc_hd__a21bo_1 _13556_ (.A1(_06265_),
    .A2(_06268_),
    .B1_N(_06266_),
    .X(_06305_));
 sky130_fd_sc_hd__and4_1 _13557_ (.A(_06195_),
    .B(\top_inst.grid_inst.data_path_wires[2][5] ),
    .C(_06202_),
    .D(_06200_),
    .X(_06306_));
 sky130_fd_sc_hd__a22oi_1 _13558_ (.A1(\top_inst.grid_inst.data_path_wires[2][5] ),
    .A2(_06202_),
    .B1(_06200_),
    .B2(_06195_),
    .Y(_06307_));
 sky130_fd_sc_hd__nor2_1 _13559_ (.A(_06306_),
    .B(_06307_),
    .Y(_06308_));
 sky130_fd_sc_hd__and2_1 _13560_ (.A(_06305_),
    .B(_06308_),
    .X(_06309_));
 sky130_fd_sc_hd__nor2_1 _13561_ (.A(_06305_),
    .B(_06308_),
    .Y(_06310_));
 sky130_fd_sc_hd__nor2_1 _13562_ (.A(_06309_),
    .B(_06310_),
    .Y(_06311_));
 sky130_fd_sc_hd__xnor2_2 _13563_ (.A(_06273_),
    .B(_06311_),
    .Y(_06312_));
 sky130_fd_sc_hd__xnor2_2 _13564_ (.A(_06304_),
    .B(_06312_),
    .Y(_06313_));
 sky130_fd_sc_hd__xor2_1 _13565_ (.A(_06293_),
    .B(_06313_),
    .X(_06314_));
 sky130_fd_sc_hd__a21oi_2 _13566_ (.A1(_06290_),
    .A2(_06291_),
    .B1(_06314_),
    .Y(_06315_));
 sky130_fd_sc_hd__and3_1 _13567_ (.A(_06290_),
    .B(_06291_),
    .C(_06314_),
    .X(_06316_));
 sky130_fd_sc_hd__inv_2 _13568_ (.A(_06278_),
    .Y(_06317_));
 sky130_fd_sc_hd__and2b_1 _13569_ (.A_N(_06280_),
    .B(_06279_),
    .X(_06318_));
 sky130_fd_sc_hd__a21oi_1 _13570_ (.A1(_06263_),
    .A2(_06317_),
    .B1(_06318_),
    .Y(_06319_));
 sky130_fd_sc_hd__nor3_2 _13571_ (.A(_06315_),
    .B(_06316_),
    .C(_06319_),
    .Y(_06320_));
 sky130_fd_sc_hd__o21a_1 _13572_ (.A1(_06315_),
    .A2(_06316_),
    .B1(_06319_),
    .X(_06321_));
 sky130_fd_sc_hd__a211oi_2 _13573_ (.A1(_06289_),
    .A2(_06285_),
    .B1(_06320_),
    .C1(_06321_),
    .Y(_06322_));
 sky130_fd_sc_hd__o211a_1 _13574_ (.A1(_06320_),
    .A2(_06321_),
    .B1(_06289_),
    .C1(_06285_),
    .X(_06323_));
 sky130_fd_sc_hd__or2_1 _13575_ (.A(_05325_),
    .B(_06323_),
    .X(_06324_));
 sky130_fd_sc_hd__a2bb2o_1 _13576_ (.A1_N(_06322_),
    .A2_N(_06324_),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[6] ),
    .B2(_05327_),
    .X(_06325_));
 sky130_fd_sc_hd__and2_1 _13577_ (.A(_05886_),
    .B(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__clkbuf_1 _13578_ (.A(_06326_),
    .X(_00373_));
 sky130_fd_sc_hd__nor2_1 _13579_ (.A(_06297_),
    .B(_06302_),
    .Y(_06327_));
 sky130_fd_sc_hd__nand2_1 _13580_ (.A(\top_inst.grid_inst.data_path_wires[2][1] ),
    .B(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[6] ),
    .Y(_06328_));
 sky130_fd_sc_hd__or2b_1 _13581_ (.A(\top_inst.grid_inst.data_path_wires[2][0] ),
    .B_N(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[7] ),
    .X(_06329_));
 sky130_fd_sc_hd__xnor2_1 _13582_ (.A(_06328_),
    .B(_06329_),
    .Y(_06330_));
 sky130_fd_sc_hd__nand2_1 _13583_ (.A(_06186_),
    .B(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[5] ),
    .Y(_06331_));
 sky130_fd_sc_hd__xnor2_1 _13584_ (.A(_06330_),
    .B(_06331_),
    .Y(_06332_));
 sky130_fd_sc_hd__xor2_1 _13585_ (.A(_06296_),
    .B(_06332_),
    .X(_06333_));
 sky130_fd_sc_hd__a22o_1 _13586_ (.A1(_06188_),
    .A2(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[2][4] ),
    .X(_06334_));
 sky130_fd_sc_hd__nand4_4 _13587_ (.A(\top_inst.grid_inst.data_path_wires[2][4] ),
    .B(_06188_),
    .C(_06210_),
    .D(_06208_),
    .Y(_06335_));
 sky130_fd_sc_hd__a22o_1 _13588_ (.A1(\top_inst.grid_inst.data_path_wires[2][5] ),
    .A2(_06205_),
    .B1(_06334_),
    .B2(_06335_),
    .X(_06336_));
 sky130_fd_sc_hd__nand4_2 _13589_ (.A(_06193_),
    .B(_06205_),
    .C(_06334_),
    .D(_06335_),
    .Y(_06337_));
 sky130_fd_sc_hd__nand2_1 _13590_ (.A(_06336_),
    .B(_06337_),
    .Y(_06338_));
 sky130_fd_sc_hd__xnor2_1 _13591_ (.A(_06333_),
    .B(_06338_),
    .Y(_06339_));
 sky130_fd_sc_hd__xnor2_1 _13592_ (.A(_06327_),
    .B(_06339_),
    .Y(_06340_));
 sky130_fd_sc_hd__nand2_1 _13593_ (.A(_06299_),
    .B(_06301_),
    .Y(_06341_));
 sky130_fd_sc_hd__a22o_1 _13594_ (.A1(\top_inst.grid_inst.data_path_wires[2][6] ),
    .A2(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[2][7] ),
    .X(_06342_));
 sky130_fd_sc_hd__and3_1 _13595_ (.A(\top_inst.grid_inst.data_path_wires[2][7] ),
    .B(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[1] ),
    .C(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[0] ),
    .X(_06343_));
 sky130_fd_sc_hd__nand2_1 _13596_ (.A(_06195_),
    .B(_06343_),
    .Y(_06344_));
 sky130_fd_sc_hd__and3_1 _13597_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[7] ),
    .B(_06342_),
    .C(_06344_),
    .X(_06345_));
 sky130_fd_sc_hd__a21oi_1 _13598_ (.A1(_06342_),
    .A2(_06344_),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[7] ),
    .Y(_06346_));
 sky130_fd_sc_hd__or2_1 _13599_ (.A(_06345_),
    .B(_06346_),
    .X(_06347_));
 sky130_fd_sc_hd__xnor2_1 _13600_ (.A(_06341_),
    .B(_06347_),
    .Y(_06348_));
 sky130_fd_sc_hd__xnor2_1 _13601_ (.A(_06306_),
    .B(_06348_),
    .Y(_06349_));
 sky130_fd_sc_hd__xor2_1 _13602_ (.A(_06340_),
    .B(_06349_),
    .X(_06350_));
 sky130_fd_sc_hd__or2_1 _13603_ (.A(_06294_),
    .B(_06303_),
    .X(_06351_));
 sky130_fd_sc_hd__o21ai_1 _13604_ (.A1(_06304_),
    .A2(_06312_),
    .B1(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__xnor2_1 _13605_ (.A(_06350_),
    .B(_06352_),
    .Y(_06353_));
 sky130_fd_sc_hd__a21o_1 _13606_ (.A1(_06273_),
    .A2(_06311_),
    .B1(_06309_),
    .X(_06354_));
 sky130_fd_sc_hd__xnor2_1 _13607_ (.A(_06353_),
    .B(_06354_),
    .Y(_06355_));
 sky130_fd_sc_hd__inv_2 _13608_ (.A(_06313_),
    .Y(_06356_));
 sky130_fd_sc_hd__a21oi_1 _13609_ (.A1(_06293_),
    .A2(_06356_),
    .B1(_06315_),
    .Y(_06357_));
 sky130_fd_sc_hd__xnor2_1 _13610_ (.A(_06355_),
    .B(_06357_),
    .Y(_06358_));
 sky130_fd_sc_hd__or3_1 _13611_ (.A(_06320_),
    .B(_06322_),
    .C(_06358_),
    .X(_06359_));
 sky130_fd_sc_hd__o21ai_2 _13612_ (.A1(_06320_),
    .A2(_06322_),
    .B1(_06358_),
    .Y(_06360_));
 sky130_fd_sc_hd__and2_1 _13613_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[7] ),
    .B(_05326_),
    .X(_06361_));
 sky130_fd_sc_hd__a31o_1 _13614_ (.A1(_05887_),
    .A2(_06359_),
    .A3(_06360_),
    .B1(_06361_),
    .X(_06362_));
 sky130_fd_sc_hd__and2_1 _13615_ (.A(_05886_),
    .B(_06362_),
    .X(_06363_));
 sky130_fd_sc_hd__clkbuf_1 _13616_ (.A(_06363_),
    .X(_00374_));
 sky130_fd_sc_hd__buf_4 _13617_ (.A(_04869_),
    .X(_06364_));
 sky130_fd_sc_hd__or2b_1 _13618_ (.A(_06357_),
    .B_N(_06355_),
    .X(_06365_));
 sky130_fd_sc_hd__and2b_1 _13619_ (.A_N(\top_inst.grid_inst.data_path_wires[2][1] ),
    .B(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[7] ),
    .X(_06366_));
 sky130_fd_sc_hd__a21oi_1 _13620_ (.A1(_06186_),
    .A2(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[6] ),
    .B1(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__and3_1 _13621_ (.A(\top_inst.grid_inst.data_path_wires[2][2] ),
    .B(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[6] ),
    .C(_06366_),
    .X(_06368_));
 sky130_fd_sc_hd__nor2_1 _13622_ (.A(_06367_),
    .B(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__nand2_1 _13623_ (.A(_06188_),
    .B(_06212_),
    .Y(_06370_));
 sky130_fd_sc_hd__xnor2_1 _13624_ (.A(_06369_),
    .B(_06370_),
    .Y(_06371_));
 sky130_fd_sc_hd__nor2_1 _13625_ (.A(_06330_),
    .B(_06331_),
    .Y(_06372_));
 sky130_fd_sc_hd__o21ba_1 _13626_ (.A1(_06328_),
    .A2(_06329_),
    .B1_N(_06372_),
    .X(_06373_));
 sky130_fd_sc_hd__xnor2_1 _13627_ (.A(_06371_),
    .B(_06373_),
    .Y(_06374_));
 sky130_fd_sc_hd__a22o_1 _13628_ (.A1(\top_inst.grid_inst.data_path_wires[2][4] ),
    .A2(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[2][5] ),
    .X(_06375_));
 sky130_fd_sc_hd__nand4_1 _13629_ (.A(\top_inst.grid_inst.data_path_wires[2][5] ),
    .B(_06190_),
    .C(_06210_),
    .D(_06208_),
    .Y(_06376_));
 sky130_fd_sc_hd__a22oi_1 _13630_ (.A1(_06195_),
    .A2(_06205_),
    .B1(_06375_),
    .B2(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__and4_1 _13631_ (.A(_06195_),
    .B(_06205_),
    .C(_06375_),
    .D(_06376_),
    .X(_06378_));
 sky130_fd_sc_hd__or2_1 _13632_ (.A(_06377_),
    .B(_06378_),
    .X(_06379_));
 sky130_fd_sc_hd__xnor2_1 _13633_ (.A(_06374_),
    .B(_06379_),
    .Y(_06380_));
 sky130_fd_sc_hd__and3_1 _13634_ (.A(_06333_),
    .B(_06336_),
    .C(_06337_),
    .X(_06381_));
 sky130_fd_sc_hd__o21ba_1 _13635_ (.A1(_06296_),
    .A2(_06332_),
    .B1_N(_06381_),
    .X(_06382_));
 sky130_fd_sc_hd__xnor2_1 _13636_ (.A(_06380_),
    .B(_06382_),
    .Y(_06383_));
 sky130_fd_sc_hd__and2_1 _13637_ (.A(_06196_),
    .B(_06343_),
    .X(_06384_));
 sky130_fd_sc_hd__o21ai_4 _13638_ (.A1(_06202_),
    .A2(_06200_),
    .B1(\top_inst.grid_inst.data_path_wires[2][7] ),
    .Y(_06385_));
 sky130_fd_sc_hd__or2_1 _13639_ (.A(_06343_),
    .B(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__a21o_1 _13640_ (.A1(_06335_),
    .A2(_06337_),
    .B1(_06386_),
    .X(_06387_));
 sky130_fd_sc_hd__nand3_1 _13641_ (.A(_06335_),
    .B(_06337_),
    .C(_06386_),
    .Y(_06388_));
 sky130_fd_sc_hd__o211a_1 _13642_ (.A1(_06384_),
    .A2(_06345_),
    .B1(_06387_),
    .C1(_06388_),
    .X(_06389_));
 sky130_fd_sc_hd__nor2_1 _13643_ (.A(_06384_),
    .B(_06345_),
    .Y(_06390_));
 sky130_fd_sc_hd__a21boi_1 _13644_ (.A1(_06387_),
    .A2(_06388_),
    .B1_N(_06390_),
    .Y(_06391_));
 sky130_fd_sc_hd__nor2_1 _13645_ (.A(_06389_),
    .B(_06391_),
    .Y(_06392_));
 sky130_fd_sc_hd__xnor2_1 _13646_ (.A(_06383_),
    .B(_06392_),
    .Y(_06393_));
 sky130_fd_sc_hd__nand2_1 _13647_ (.A(_06327_),
    .B(_06339_),
    .Y(_06394_));
 sky130_fd_sc_hd__o21a_1 _13648_ (.A1(_06340_),
    .A2(_06349_),
    .B1(_06394_),
    .X(_06395_));
 sky130_fd_sc_hd__xnor2_1 _13649_ (.A(_06393_),
    .B(_06395_),
    .Y(_06396_));
 sky130_fd_sc_hd__or2b_1 _13650_ (.A(_06347_),
    .B_N(_06341_),
    .X(_06397_));
 sky130_fd_sc_hd__a21boi_1 _13651_ (.A1(_06306_),
    .A2(_06348_),
    .B1_N(_06397_),
    .Y(_06398_));
 sky130_fd_sc_hd__xnor2_1 _13652_ (.A(_06396_),
    .B(_06398_),
    .Y(_06399_));
 sky130_fd_sc_hd__or2b_1 _13653_ (.A(_06353_),
    .B_N(_06354_),
    .X(_06400_));
 sky130_fd_sc_hd__a21boi_1 _13654_ (.A1(_06350_),
    .A2(_06352_),
    .B1_N(_06400_),
    .Y(_06401_));
 sky130_fd_sc_hd__xnor2_1 _13655_ (.A(_06399_),
    .B(_06401_),
    .Y(_06402_));
 sky130_fd_sc_hd__a21o_1 _13656_ (.A1(_06365_),
    .A2(_06360_),
    .B1(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__clkbuf_8 _13657_ (.A(_05325_),
    .X(_06404_));
 sky130_fd_sc_hd__a31oi_1 _13658_ (.A1(_06365_),
    .A2(_06360_),
    .A3(_06402_),
    .B1(_06404_),
    .Y(_06405_));
 sky130_fd_sc_hd__a22o_1 _13659_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[8] ),
    .A2(_06242_),
    .B1(_06403_),
    .B2(_06405_),
    .X(_06406_));
 sky130_fd_sc_hd__and2_1 _13660_ (.A(_06364_),
    .B(_06406_),
    .X(_06407_));
 sky130_fd_sc_hd__clkbuf_1 _13661_ (.A(_06407_),
    .X(_00375_));
 sky130_fd_sc_hd__nor2_1 _13662_ (.A(_06399_),
    .B(_06401_),
    .Y(_06408_));
 sky130_fd_sc_hd__inv_2 _13663_ (.A(_06408_),
    .Y(_06409_));
 sky130_fd_sc_hd__and2b_1 _13664_ (.A_N(\top_inst.grid_inst.data_path_wires[2][2] ),
    .B(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[7] ),
    .X(_06410_));
 sky130_fd_sc_hd__a21oi_1 _13665_ (.A1(_06188_),
    .A2(_06214_),
    .B1(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__and3_1 _13666_ (.A(_06188_),
    .B(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[6] ),
    .C(_06410_),
    .X(_06412_));
 sky130_fd_sc_hd__nor2_1 _13667_ (.A(_06411_),
    .B(_06412_),
    .Y(_06413_));
 sky130_fd_sc_hd__nand2_1 _13668_ (.A(_06190_),
    .B(_06212_),
    .Y(_06414_));
 sky130_fd_sc_hd__xnor2_1 _13669_ (.A(_06413_),
    .B(_06414_),
    .Y(_06415_));
 sky130_fd_sc_hd__o21ba_1 _13670_ (.A1(_06367_),
    .A2(_06370_),
    .B1_N(_06368_),
    .X(_06416_));
 sky130_fd_sc_hd__xor2_1 _13671_ (.A(_06415_),
    .B(_06416_),
    .X(_06417_));
 sky130_fd_sc_hd__a22oi_2 _13672_ (.A1(_06193_),
    .A2(_06210_),
    .B1(_06208_),
    .B2(_06195_),
    .Y(_06418_));
 sky130_fd_sc_hd__and4_1 _13673_ (.A(_06195_),
    .B(\top_inst.grid_inst.data_path_wires[2][5] ),
    .C(_06210_),
    .D(_06208_),
    .X(_06419_));
 sky130_fd_sc_hd__nor2_1 _13674_ (.A(_06418_),
    .B(_06419_),
    .Y(_06420_));
 sky130_fd_sc_hd__nand2_2 _13675_ (.A(_06198_),
    .B(_06205_),
    .Y(_06421_));
 sky130_fd_sc_hd__xor2_1 _13676_ (.A(_06420_),
    .B(_06421_),
    .X(_06422_));
 sky130_fd_sc_hd__xor2_1 _13677_ (.A(_06417_),
    .B(_06422_),
    .X(_06423_));
 sky130_fd_sc_hd__inv_2 _13678_ (.A(_06373_),
    .Y(_06424_));
 sky130_fd_sc_hd__or3b_1 _13679_ (.A(_06377_),
    .B(_06378_),
    .C_N(_06374_),
    .X(_06425_));
 sky130_fd_sc_hd__a21boi_1 _13680_ (.A1(_06371_),
    .A2(_06424_),
    .B1_N(_06425_),
    .Y(_06426_));
 sky130_fd_sc_hd__xnor2_1 _13681_ (.A(_06423_),
    .B(_06426_),
    .Y(_06427_));
 sky130_fd_sc_hd__and4_1 _13682_ (.A(_06193_),
    .B(_06190_),
    .C(_06210_),
    .D(_06208_),
    .X(_06428_));
 sky130_fd_sc_hd__nor2_1 _13683_ (.A(_06428_),
    .B(_06378_),
    .Y(_06429_));
 sky130_fd_sc_hd__nor2_1 _13684_ (.A(_06385_),
    .B(_06429_),
    .Y(_06430_));
 sky130_fd_sc_hd__and2_1 _13685_ (.A(_06385_),
    .B(_06429_),
    .X(_06431_));
 sky130_fd_sc_hd__nor2_1 _13686_ (.A(_06430_),
    .B(_06431_),
    .Y(_06432_));
 sky130_fd_sc_hd__xnor2_1 _13687_ (.A(_06427_),
    .B(_06432_),
    .Y(_06433_));
 sky130_fd_sc_hd__and2b_1 _13688_ (.A_N(_06382_),
    .B(_06380_),
    .X(_06434_));
 sky130_fd_sc_hd__a21oi_1 _13689_ (.A1(_06383_),
    .A2(_06392_),
    .B1(_06434_),
    .Y(_06435_));
 sky130_fd_sc_hd__xnor2_1 _13690_ (.A(_06433_),
    .B(_06435_),
    .Y(_06436_));
 sky130_fd_sc_hd__and3_1 _13691_ (.A(_06335_),
    .B(_06337_),
    .C(_06386_),
    .X(_06437_));
 sky130_fd_sc_hd__o21a_1 _13692_ (.A1(_06390_),
    .A2(_06437_),
    .B1(_06387_),
    .X(_06438_));
 sky130_fd_sc_hd__xnor2_1 _13693_ (.A(_06436_),
    .B(_06438_),
    .Y(_06439_));
 sky130_fd_sc_hd__or2_1 _13694_ (.A(_06393_),
    .B(_06395_),
    .X(_06440_));
 sky130_fd_sc_hd__o21a_1 _13695_ (.A1(_06396_),
    .A2(_06398_),
    .B1(_06440_),
    .X(_06441_));
 sky130_fd_sc_hd__xnor2_1 _13696_ (.A(_06439_),
    .B(_06441_),
    .Y(_06442_));
 sky130_fd_sc_hd__a21o_1 _13697_ (.A1(_06409_),
    .A2(_06403_),
    .B1(_06442_),
    .X(_06443_));
 sky130_fd_sc_hd__nand3_1 _13698_ (.A(_06409_),
    .B(_06403_),
    .C(_06442_),
    .Y(_06444_));
 sky130_fd_sc_hd__a21o_1 _13699_ (.A1(_06443_),
    .A2(_06444_),
    .B1(_05328_),
    .X(_06445_));
 sky130_fd_sc_hd__clkbuf_4 _13700_ (.A(_05260_),
    .X(_06446_));
 sky130_fd_sc_hd__o211a_1 _13701_ (.A1(net1061),
    .A2(_05788_),
    .B1(_06445_),
    .C1(_06446_),
    .X(_00376_));
 sky130_fd_sc_hd__or2_1 _13702_ (.A(_06439_),
    .B(_06441_),
    .X(_06447_));
 sky130_fd_sc_hd__or2b_1 _13703_ (.A(_06416_),
    .B_N(_06415_),
    .X(_06448_));
 sky130_fd_sc_hd__o21a_1 _13704_ (.A1(_06417_),
    .A2(_06422_),
    .B1(_06448_),
    .X(_06449_));
 sky130_fd_sc_hd__and2b_1 _13705_ (.A_N(\top_inst.grid_inst.data_path_wires[2][3] ),
    .B(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[7] ),
    .X(_06450_));
 sky130_fd_sc_hd__a21oi_1 _13706_ (.A1(_06190_),
    .A2(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[6] ),
    .B1(_06450_),
    .Y(_06451_));
 sky130_fd_sc_hd__and3_1 _13707_ (.A(\top_inst.grid_inst.data_path_wires[2][4] ),
    .B(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[6] ),
    .C(_06450_),
    .X(_06452_));
 sky130_fd_sc_hd__nor2_1 _13708_ (.A(_06451_),
    .B(_06452_),
    .Y(_06453_));
 sky130_fd_sc_hd__nand2_1 _13709_ (.A(\top_inst.grid_inst.data_path_wires[2][5] ),
    .B(_06212_),
    .Y(_06454_));
 sky130_fd_sc_hd__xnor2_1 _13710_ (.A(_06453_),
    .B(_06454_),
    .Y(_06455_));
 sky130_fd_sc_hd__o21ba_1 _13711_ (.A1(_06411_),
    .A2(_06414_),
    .B1_N(_06412_),
    .X(_06456_));
 sky130_fd_sc_hd__xor2_1 _13712_ (.A(_06455_),
    .B(_06456_),
    .X(_06457_));
 sky130_fd_sc_hd__and3_2 _13713_ (.A(\top_inst.grid_inst.data_path_wires[2][7] ),
    .B(_06210_),
    .C(_06208_),
    .X(_06458_));
 sky130_fd_sc_hd__a22oi_1 _13714_ (.A1(_06195_),
    .A2(_06210_),
    .B1(_06208_),
    .B2(\top_inst.grid_inst.data_path_wires[2][7] ),
    .Y(_06459_));
 sky130_fd_sc_hd__a21oi_1 _13715_ (.A1(_06196_),
    .A2(_06458_),
    .B1(_06459_),
    .Y(_06460_));
 sky130_fd_sc_hd__xnor2_1 _13716_ (.A(_06421_),
    .B(_06460_),
    .Y(_06461_));
 sky130_fd_sc_hd__xnor2_1 _13717_ (.A(_06457_),
    .B(_06461_),
    .Y(_06462_));
 sky130_fd_sc_hd__and2b_1 _13718_ (.A_N(_06449_),
    .B(_06462_),
    .X(_06463_));
 sky130_fd_sc_hd__and2b_1 _13719_ (.A_N(_06462_),
    .B(_06449_),
    .X(_06464_));
 sky130_fd_sc_hd__nor2_1 _13720_ (.A(_06463_),
    .B(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__o21ba_1 _13721_ (.A1(_06418_),
    .A2(_06421_),
    .B1_N(_06419_),
    .X(_06466_));
 sky130_fd_sc_hd__nor2_1 _13722_ (.A(_06385_),
    .B(_06466_),
    .Y(_06467_));
 sky130_fd_sc_hd__and2_1 _13723_ (.A(_06385_),
    .B(_06466_),
    .X(_06468_));
 sky130_fd_sc_hd__nor2_1 _13724_ (.A(_06467_),
    .B(_06468_),
    .Y(_06469_));
 sky130_fd_sc_hd__xnor2_1 _13725_ (.A(_06465_),
    .B(_06469_),
    .Y(_06470_));
 sky130_fd_sc_hd__and2b_1 _13726_ (.A_N(_06426_),
    .B(_06423_),
    .X(_06471_));
 sky130_fd_sc_hd__a21oi_1 _13727_ (.A1(_06427_),
    .A2(_06432_),
    .B1(_06471_),
    .Y(_06472_));
 sky130_fd_sc_hd__xor2_1 _13728_ (.A(_06470_),
    .B(_06472_),
    .X(_06473_));
 sky130_fd_sc_hd__xnor2_1 _13729_ (.A(_06430_),
    .B(_06473_),
    .Y(_06474_));
 sky130_fd_sc_hd__or2_1 _13730_ (.A(_06433_),
    .B(_06435_),
    .X(_06475_));
 sky130_fd_sc_hd__o21a_1 _13731_ (.A1(_06436_),
    .A2(_06438_),
    .B1(_06475_),
    .X(_06476_));
 sky130_fd_sc_hd__nor2_1 _13732_ (.A(_06474_),
    .B(_06476_),
    .Y(_06477_));
 sky130_fd_sc_hd__and2_1 _13733_ (.A(_06474_),
    .B(_06476_),
    .X(_06478_));
 sky130_fd_sc_hd__or2_1 _13734_ (.A(_06477_),
    .B(_06478_),
    .X(_06479_));
 sky130_fd_sc_hd__a21o_1 _13735_ (.A1(_06447_),
    .A2(_06443_),
    .B1(_06479_),
    .X(_06480_));
 sky130_fd_sc_hd__a31oi_1 _13736_ (.A1(_06447_),
    .A2(_06443_),
    .A3(_06479_),
    .B1(_06404_),
    .Y(_06481_));
 sky130_fd_sc_hd__a22o_1 _13737_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[10] ),
    .A2(_06242_),
    .B1(_06480_),
    .B2(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__and2_1 _13738_ (.A(_06364_),
    .B(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__clkbuf_1 _13739_ (.A(_06483_),
    .X(_00377_));
 sky130_fd_sc_hd__inv_2 _13740_ (.A(_06477_),
    .Y(_06484_));
 sky130_fd_sc_hd__and2b_1 _13741_ (.A_N(\top_inst.grid_inst.data_path_wires[2][4] ),
    .B(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[7] ),
    .X(_06485_));
 sky130_fd_sc_hd__a21oi_1 _13742_ (.A1(_06193_),
    .A2(_06214_),
    .B1(_06485_),
    .Y(_06486_));
 sky130_fd_sc_hd__and3_1 _13743_ (.A(_06193_),
    .B(_06214_),
    .C(_06485_),
    .X(_06487_));
 sky130_fd_sc_hd__nor2_1 _13744_ (.A(_06486_),
    .B(_06487_),
    .Y(_06488_));
 sky130_fd_sc_hd__nand2_1 _13745_ (.A(_06196_),
    .B(_06212_),
    .Y(_06489_));
 sky130_fd_sc_hd__xnor2_1 _13746_ (.A(_06488_),
    .B(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__o21ba_1 _13747_ (.A1(_06451_),
    .A2(_06454_),
    .B1_N(_06452_),
    .X(_06491_));
 sky130_fd_sc_hd__xnor2_1 _13748_ (.A(_06490_),
    .B(_06491_),
    .Y(_06492_));
 sky130_fd_sc_hd__o21ai_1 _13749_ (.A1(_06210_),
    .A2(_06208_),
    .B1(_06198_),
    .Y(_06493_));
 sky130_fd_sc_hd__nor3_1 _13750_ (.A(_06421_),
    .B(_06458_),
    .C(_06493_),
    .Y(_06494_));
 sky130_fd_sc_hd__o21a_1 _13751_ (.A1(_06458_),
    .A2(_06493_),
    .B1(_06421_),
    .X(_06495_));
 sky130_fd_sc_hd__nor2_2 _13752_ (.A(_06494_),
    .B(_06495_),
    .Y(_06496_));
 sky130_fd_sc_hd__or2_1 _13753_ (.A(_06492_),
    .B(_06496_),
    .X(_06497_));
 sky130_fd_sc_hd__nand2_1 _13754_ (.A(_06492_),
    .B(_06496_),
    .Y(_06498_));
 sky130_fd_sc_hd__nand2_1 _13755_ (.A(_06497_),
    .B(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__or2b_1 _13756_ (.A(_06455_),
    .B_N(_06456_),
    .X(_06500_));
 sky130_fd_sc_hd__and2b_1 _13757_ (.A_N(_06456_),
    .B(_06455_),
    .X(_06501_));
 sky130_fd_sc_hd__a21oi_1 _13758_ (.A1(_06500_),
    .A2(_06461_),
    .B1(_06501_),
    .Y(_06502_));
 sky130_fd_sc_hd__nor2_1 _13759_ (.A(_06499_),
    .B(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__and2_1 _13760_ (.A(_06499_),
    .B(_06502_),
    .X(_06504_));
 sky130_fd_sc_hd__nor2_1 _13761_ (.A(_06503_),
    .B(_06504_),
    .Y(_06505_));
 sky130_fd_sc_hd__o2bb2a_1 _13762_ (.A1_N(_06196_),
    .A2_N(_06458_),
    .B1(_06459_),
    .B2(_06421_),
    .X(_06506_));
 sky130_fd_sc_hd__nor2_1 _13763_ (.A(_06385_),
    .B(_06506_),
    .Y(_06507_));
 sky130_fd_sc_hd__and2_1 _13764_ (.A(_06385_),
    .B(_06506_),
    .X(_06508_));
 sky130_fd_sc_hd__nor2_1 _13765_ (.A(_06507_),
    .B(_06508_),
    .Y(_06509_));
 sky130_fd_sc_hd__xnor2_1 _13766_ (.A(_06505_),
    .B(_06509_),
    .Y(_06510_));
 sky130_fd_sc_hd__a21oi_1 _13767_ (.A1(_06465_),
    .A2(_06469_),
    .B1(_06463_),
    .Y(_06511_));
 sky130_fd_sc_hd__nor2_1 _13768_ (.A(_06510_),
    .B(_06511_),
    .Y(_06512_));
 sky130_fd_sc_hd__and2_1 _13769_ (.A(_06510_),
    .B(_06511_),
    .X(_06513_));
 sky130_fd_sc_hd__nor2_1 _13770_ (.A(_06512_),
    .B(_06513_),
    .Y(_06514_));
 sky130_fd_sc_hd__xnor2_1 _13771_ (.A(_06467_),
    .B(_06514_),
    .Y(_06515_));
 sky130_fd_sc_hd__nor2_1 _13772_ (.A(_06470_),
    .B(_06472_),
    .Y(_06516_));
 sky130_fd_sc_hd__a21oi_1 _13773_ (.A1(_06430_),
    .A2(_06473_),
    .B1(_06516_),
    .Y(_06517_));
 sky130_fd_sc_hd__xnor2_1 _13774_ (.A(_06515_),
    .B(_06517_),
    .Y(_06518_));
 sky130_fd_sc_hd__a21o_1 _13775_ (.A1(_06484_),
    .A2(_06480_),
    .B1(_06518_),
    .X(_06519_));
 sky130_fd_sc_hd__nand3_1 _13776_ (.A(_06484_),
    .B(_06480_),
    .C(_06518_),
    .Y(_06520_));
 sky130_fd_sc_hd__a21o_1 _13777_ (.A1(_06519_),
    .A2(_06520_),
    .B1(_05328_),
    .X(_06521_));
 sky130_fd_sc_hd__o211a_1 _13778_ (.A1(net1052),
    .A2(_05788_),
    .B1(_06521_),
    .C1(_06446_),
    .X(_00378_));
 sky130_fd_sc_hd__or2_1 _13779_ (.A(_06515_),
    .B(_06517_),
    .X(_06522_));
 sky130_fd_sc_hd__or2b_1 _13780_ (.A(_06491_),
    .B_N(_06490_),
    .X(_06523_));
 sky130_fd_sc_hd__inv_2 _13781_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[7] ),
    .Y(_06524_));
 sky130_fd_sc_hd__o2bb2a_1 _13782_ (.A1_N(_06196_),
    .A2_N(_06214_),
    .B1(_06524_),
    .B2(_06193_),
    .X(_06525_));
 sky130_fd_sc_hd__and4b_1 _13783_ (.A_N(_06193_),
    .B(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[7] ),
    .C(_06214_),
    .D(_06195_),
    .X(_06526_));
 sky130_fd_sc_hd__nand2_1 _13784_ (.A(_06198_),
    .B(_06212_),
    .Y(_06527_));
 sky130_fd_sc_hd__o21a_1 _13785_ (.A1(_06525_),
    .A2(_06526_),
    .B1(_06527_),
    .X(_06528_));
 sky130_fd_sc_hd__nor2_1 _13786_ (.A(_06525_),
    .B(_06526_),
    .Y(_06529_));
 sky130_fd_sc_hd__and3_1 _13787_ (.A(_06198_),
    .B(_06212_),
    .C(_06529_),
    .X(_06530_));
 sky130_fd_sc_hd__nor2_1 _13788_ (.A(_06528_),
    .B(_06530_),
    .Y(_06531_));
 sky130_fd_sc_hd__o21ba_1 _13789_ (.A1(_06486_),
    .A2(_06489_),
    .B1_N(_06487_),
    .X(_06532_));
 sky130_fd_sc_hd__xnor2_1 _13790_ (.A(_06531_),
    .B(_06532_),
    .Y(_06533_));
 sky130_fd_sc_hd__xnor2_1 _13791_ (.A(_06496_),
    .B(_06533_),
    .Y(_06534_));
 sky130_fd_sc_hd__a21o_1 _13792_ (.A1(_06523_),
    .A2(_06498_),
    .B1(_06534_),
    .X(_06535_));
 sky130_fd_sc_hd__nand3_1 _13793_ (.A(_06523_),
    .B(_06498_),
    .C(_06534_),
    .Y(_06536_));
 sky130_fd_sc_hd__nand2_1 _13794_ (.A(_06535_),
    .B(_06536_),
    .Y(_06537_));
 sky130_fd_sc_hd__o21a_1 _13795_ (.A1(_06202_),
    .A2(_06200_),
    .B1(_06198_),
    .X(_06538_));
 sky130_fd_sc_hd__o21ai_2 _13796_ (.A1(_06458_),
    .A2(net181),
    .B1(_06538_),
    .Y(_06539_));
 sky130_fd_sc_hd__or3_2 _13797_ (.A(_06538_),
    .B(_06458_),
    .C(net181),
    .X(_06540_));
 sky130_fd_sc_hd__nand2_2 _13798_ (.A(_06539_),
    .B(_06540_),
    .Y(_06541_));
 sky130_fd_sc_hd__inv_2 _13799_ (.A(_06541_),
    .Y(_06542_));
 sky130_fd_sc_hd__xnor2_1 _13800_ (.A(_06537_),
    .B(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__a21oi_1 _13801_ (.A1(_06505_),
    .A2(_06509_),
    .B1(_06503_),
    .Y(_06544_));
 sky130_fd_sc_hd__xnor2_1 _13802_ (.A(_06543_),
    .B(_06544_),
    .Y(_06545_));
 sky130_fd_sc_hd__xnor2_1 _13803_ (.A(_06507_),
    .B(_06545_),
    .Y(_06546_));
 sky130_fd_sc_hd__a21oi_1 _13804_ (.A1(_06467_),
    .A2(_06514_),
    .B1(_06512_),
    .Y(_06547_));
 sky130_fd_sc_hd__or2_1 _13805_ (.A(_06546_),
    .B(_06547_),
    .X(_06548_));
 sky130_fd_sc_hd__nand2_1 _13806_ (.A(_06546_),
    .B(_06547_),
    .Y(_06549_));
 sky130_fd_sc_hd__nand2_1 _13807_ (.A(_06548_),
    .B(_06549_),
    .Y(_06550_));
 sky130_fd_sc_hd__a21o_1 _13808_ (.A1(_06522_),
    .A2(_06519_),
    .B1(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__a31oi_1 _13809_ (.A1(_06522_),
    .A2(_06519_),
    .A3(_06550_),
    .B1(_06404_),
    .Y(_06552_));
 sky130_fd_sc_hd__a22o_1 _13810_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[12] ),
    .A2(_06242_),
    .B1(_06551_),
    .B2(_06552_),
    .X(_06553_));
 sky130_fd_sc_hd__and2_1 _13811_ (.A(_06364_),
    .B(_06553_),
    .X(_06554_));
 sky130_fd_sc_hd__clkbuf_1 _13812_ (.A(_06554_),
    .X(_00379_));
 sky130_fd_sc_hd__inv_2 _13813_ (.A(_06539_),
    .Y(_06555_));
 sky130_fd_sc_hd__o21a_1 _13814_ (.A1(_06537_),
    .A2(_06541_),
    .B1(_06535_),
    .X(_06556_));
 sky130_fd_sc_hd__nand2_1 _13815_ (.A(\top_inst.grid_inst.data_path_wires[2][7] ),
    .B(_06214_),
    .Y(_06557_));
 sky130_fd_sc_hd__o21a_1 _13816_ (.A1(_06196_),
    .A2(_06524_),
    .B1(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__nor3_1 _13817_ (.A(_06196_),
    .B(_06524_),
    .C(_06557_),
    .Y(_06559_));
 sky130_fd_sc_hd__nor2_1 _13818_ (.A(_06558_),
    .B(_06559_),
    .Y(_06560_));
 sky130_fd_sc_hd__xnor2_1 _13819_ (.A(_06527_),
    .B(_06560_),
    .Y(_06561_));
 sky130_fd_sc_hd__o21ai_1 _13820_ (.A1(_06526_),
    .A2(_06530_),
    .B1(_06561_),
    .Y(_06562_));
 sky130_fd_sc_hd__or3_1 _13821_ (.A(_06526_),
    .B(_06530_),
    .C(_06561_),
    .X(_06563_));
 sky130_fd_sc_hd__and2_1 _13822_ (.A(_06562_),
    .B(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__nand2_1 _13823_ (.A(_06496_),
    .B(_06564_),
    .Y(_06565_));
 sky130_fd_sc_hd__or2_1 _13824_ (.A(_06496_),
    .B(_06564_),
    .X(_06566_));
 sky130_fd_sc_hd__nand2_1 _13825_ (.A(_06565_),
    .B(_06566_),
    .Y(_06567_));
 sky130_fd_sc_hd__or2b_1 _13826_ (.A(_06532_),
    .B_N(_06531_),
    .X(_06568_));
 sky130_fd_sc_hd__a21bo_1 _13827_ (.A1(_06496_),
    .A2(_06533_),
    .B1_N(_06568_),
    .X(_06569_));
 sky130_fd_sc_hd__xor2_1 _13828_ (.A(_06567_),
    .B(_06569_),
    .X(_06570_));
 sky130_fd_sc_hd__xnor2_1 _13829_ (.A(_06542_),
    .B(_06570_),
    .Y(_06571_));
 sky130_fd_sc_hd__and2b_1 _13830_ (.A_N(_06556_),
    .B(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__and2b_1 _13831_ (.A_N(_06571_),
    .B(_06556_),
    .X(_06573_));
 sky130_fd_sc_hd__nor2_1 _13832_ (.A(_06572_),
    .B(_06573_),
    .Y(_06574_));
 sky130_fd_sc_hd__xnor2_1 _13833_ (.A(_06555_),
    .B(_06574_),
    .Y(_06575_));
 sky130_fd_sc_hd__and2b_1 _13834_ (.A_N(_06544_),
    .B(_06543_),
    .X(_06576_));
 sky130_fd_sc_hd__a21oi_1 _13835_ (.A1(_06507_),
    .A2(_06545_),
    .B1(_06576_),
    .Y(_06577_));
 sky130_fd_sc_hd__or2_1 _13836_ (.A(_06575_),
    .B(_06577_),
    .X(_06578_));
 sky130_fd_sc_hd__nand2_1 _13837_ (.A(_06575_),
    .B(_06577_),
    .Y(_06579_));
 sky130_fd_sc_hd__nand2_1 _13838_ (.A(_06578_),
    .B(_06579_),
    .Y(_06580_));
 sky130_fd_sc_hd__and3_1 _13839_ (.A(_06548_),
    .B(_06551_),
    .C(_06580_),
    .X(_06581_));
 sky130_fd_sc_hd__a21o_1 _13840_ (.A1(_06548_),
    .A2(_06551_),
    .B1(_06580_),
    .X(_06582_));
 sky130_fd_sc_hd__nand2_1 _13841_ (.A(_06140_),
    .B(_06582_),
    .Y(_06583_));
 sky130_fd_sc_hd__a2bb2o_1 _13842_ (.A1_N(_06581_),
    .A2_N(_06583_),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[13] ),
    .B2(_05327_),
    .X(_06584_));
 sky130_fd_sc_hd__and2_1 _13843_ (.A(_06364_),
    .B(_06584_),
    .X(_06585_));
 sky130_fd_sc_hd__clkbuf_1 _13844_ (.A(_06585_),
    .X(_00380_));
 sky130_fd_sc_hd__or2b_1 _13845_ (.A(_06567_),
    .B_N(_06569_),
    .X(_06586_));
 sky130_fd_sc_hd__o21a_1 _13846_ (.A1(_06541_),
    .A2(_06570_),
    .B1(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__and3_1 _13847_ (.A(_06198_),
    .B(_06214_),
    .C(_06212_),
    .X(_06588_));
 sky130_fd_sc_hd__o21ba_1 _13848_ (.A1(_06527_),
    .A2(_06558_),
    .B1_N(_06559_),
    .X(_06589_));
 sky130_fd_sc_hd__o211a_1 _13849_ (.A1(_06198_),
    .A2(_06524_),
    .B1(_06527_),
    .C1(_06557_),
    .X(_06590_));
 sky130_fd_sc_hd__o21ba_1 _13850_ (.A1(_06588_),
    .A2(_06589_),
    .B1_N(_06590_),
    .X(_06591_));
 sky130_fd_sc_hd__xnor2_1 _13851_ (.A(_06496_),
    .B(_06591_),
    .Y(_06592_));
 sky130_fd_sc_hd__a21oi_1 _13852_ (.A1(_06562_),
    .A2(_06565_),
    .B1(_06592_),
    .Y(_06593_));
 sky130_fd_sc_hd__and3_1 _13853_ (.A(_06562_),
    .B(_06565_),
    .C(_06592_),
    .X(_06594_));
 sky130_fd_sc_hd__nor2_1 _13854_ (.A(_06593_),
    .B(_06594_),
    .Y(_06595_));
 sky130_fd_sc_hd__xnor2_1 _13855_ (.A(_06541_),
    .B(_06595_),
    .Y(_06596_));
 sky130_fd_sc_hd__and2b_1 _13856_ (.A_N(_06587_),
    .B(_06596_),
    .X(_06597_));
 sky130_fd_sc_hd__and2b_1 _13857_ (.A_N(_06596_),
    .B(_06587_),
    .X(_06598_));
 sky130_fd_sc_hd__nor2_1 _13858_ (.A(_06597_),
    .B(_06598_),
    .Y(_06599_));
 sky130_fd_sc_hd__xnor2_1 _13859_ (.A(_06555_),
    .B(_06599_),
    .Y(_06600_));
 sky130_fd_sc_hd__a21oi_1 _13860_ (.A1(_06555_),
    .A2(_06574_),
    .B1(_06572_),
    .Y(_06601_));
 sky130_fd_sc_hd__or2_1 _13861_ (.A(_06600_),
    .B(_06601_),
    .X(_06602_));
 sky130_fd_sc_hd__nand2_1 _13862_ (.A(_06600_),
    .B(_06601_),
    .Y(_06603_));
 sky130_fd_sc_hd__nand2_1 _13863_ (.A(_06602_),
    .B(_06603_),
    .Y(_06604_));
 sky130_fd_sc_hd__a21o_1 _13864_ (.A1(_06578_),
    .A2(_06582_),
    .B1(_06604_),
    .X(_06605_));
 sky130_fd_sc_hd__a31oi_1 _13865_ (.A1(_06578_),
    .A2(_06582_),
    .A3(_06604_),
    .B1(_06404_),
    .Y(_06606_));
 sky130_fd_sc_hd__a22o_1 _13866_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[14] ),
    .A2(_06242_),
    .B1(_06605_),
    .B2(_06606_),
    .X(_06607_));
 sky130_fd_sc_hd__and2_1 _13867_ (.A(_06364_),
    .B(_06607_),
    .X(_06608_));
 sky130_fd_sc_hd__clkbuf_1 _13868_ (.A(_06608_),
    .X(_00381_));
 sky130_fd_sc_hd__and3_1 _13869_ (.A(_06540_),
    .B(_06602_),
    .C(_06605_),
    .X(_06609_));
 sky130_fd_sc_hd__a21oi_1 _13870_ (.A1(_06602_),
    .A2(_06605_),
    .B1(_06540_),
    .Y(_06610_));
 sky130_fd_sc_hd__nor2_1 _13871_ (.A(_06496_),
    .B(_06591_),
    .Y(_06611_));
 sky130_fd_sc_hd__a21oi_1 _13872_ (.A1(_06555_),
    .A2(_06599_),
    .B1(_06597_),
    .Y(_06612_));
 sky130_fd_sc_hd__a21oi_1 _13873_ (.A1(_06542_),
    .A2(_06595_),
    .B1(_06593_),
    .Y(_06613_));
 sky130_fd_sc_hd__xnor2_1 _13874_ (.A(_06612_),
    .B(_06613_),
    .Y(_06614_));
 sky130_fd_sc_hd__xnor2_1 _13875_ (.A(_06611_),
    .B(_06614_),
    .Y(_06615_));
 sky130_fd_sc_hd__o21a_1 _13876_ (.A1(_06609_),
    .A2(_06610_),
    .B1(_06615_),
    .X(_06616_));
 sky130_fd_sc_hd__o31ai_1 _13877_ (.A1(_06609_),
    .A2(_06610_),
    .A3(_06615_),
    .B1(_05313_),
    .Y(_06617_));
 sky130_fd_sc_hd__o221a_1 _13878_ (.A1(net1074),
    .A2(_06169_),
    .B1(_06616_),
    .B2(_06617_),
    .C1(_06180_),
    .X(_00382_));
 sky130_fd_sc_hd__buf_2 _13879_ (.A(\top_inst.grid_inst.data_path_wires[3][0] ),
    .X(_06618_));
 sky130_fd_sc_hd__buf_6 _13880_ (.A(_04862_),
    .X(_06619_));
 sky130_fd_sc_hd__buf_2 _13881_ (.A(_06619_),
    .X(_06620_));
 sky130_fd_sc_hd__or2_1 _13882_ (.A(_06618_),
    .B(_06620_),
    .X(_06621_));
 sky130_fd_sc_hd__o211a_1 _13883_ (.A1(_06181_),
    .A2(_06192_),
    .B1(_06621_),
    .C1(_06446_),
    .X(_00383_));
 sky130_fd_sc_hd__clkbuf_4 _13884_ (.A(\top_inst.grid_inst.data_path_wires[3][1] ),
    .X(_06622_));
 sky130_fd_sc_hd__or2_1 _13885_ (.A(_06622_),
    .B(_06620_),
    .X(_06623_));
 sky130_fd_sc_hd__o211a_1 _13886_ (.A1(_06184_),
    .A2(_06192_),
    .B1(_06623_),
    .C1(_06446_),
    .X(_00384_));
 sky130_fd_sc_hd__clkbuf_4 _13887_ (.A(\top_inst.grid_inst.data_path_wires[3][2] ),
    .X(_06624_));
 sky130_fd_sc_hd__or2_1 _13888_ (.A(_06624_),
    .B(_06620_),
    .X(_06625_));
 sky130_fd_sc_hd__o211a_1 _13889_ (.A1(_06186_),
    .A2(_06192_),
    .B1(_06625_),
    .C1(_06446_),
    .X(_00385_));
 sky130_fd_sc_hd__clkbuf_4 _13890_ (.A(\top_inst.grid_inst.data_path_wires[3][3] ),
    .X(_06626_));
 sky130_fd_sc_hd__or2_1 _13891_ (.A(_06626_),
    .B(_06620_),
    .X(_06627_));
 sky130_fd_sc_hd__o211a_1 _13892_ (.A1(_06188_),
    .A2(_06192_),
    .B1(_06627_),
    .C1(_06446_),
    .X(_00386_));
 sky130_fd_sc_hd__clkbuf_4 _13893_ (.A(\top_inst.grid_inst.data_path_wires[3][4] ),
    .X(_06628_));
 sky130_fd_sc_hd__or2_1 _13894_ (.A(_06628_),
    .B(_06620_),
    .X(_06629_));
 sky130_fd_sc_hd__o211a_1 _13895_ (.A1(_06190_),
    .A2(_06192_),
    .B1(_06629_),
    .C1(_06446_),
    .X(_00387_));
 sky130_fd_sc_hd__clkbuf_4 _13896_ (.A(\top_inst.grid_inst.data_path_wires[3][5] ),
    .X(_06630_));
 sky130_fd_sc_hd__or2_1 _13897_ (.A(_06630_),
    .B(_06620_),
    .X(_06631_));
 sky130_fd_sc_hd__o211a_1 _13898_ (.A1(_06193_),
    .A2(_06192_),
    .B1(_06631_),
    .C1(_06446_),
    .X(_00388_));
 sky130_fd_sc_hd__clkbuf_4 _13899_ (.A(\top_inst.grid_inst.data_path_wires[3][6] ),
    .X(_06632_));
 sky130_fd_sc_hd__or2_1 _13900_ (.A(_06632_),
    .B(_06620_),
    .X(_06633_));
 sky130_fd_sc_hd__o211a_1 _13901_ (.A1(_06196_),
    .A2(_06192_),
    .B1(_06633_),
    .C1(_06446_),
    .X(_00389_));
 sky130_fd_sc_hd__clkbuf_4 _13902_ (.A(_05177_),
    .X(_06634_));
 sky130_fd_sc_hd__clkbuf_4 _13903_ (.A(\top_inst.grid_inst.data_path_wires[3][7] ),
    .X(_06635_));
 sky130_fd_sc_hd__or2_1 _13904_ (.A(_06635_),
    .B(_06620_),
    .X(_06636_));
 sky130_fd_sc_hd__o211a_1 _13905_ (.A1(_06198_),
    .A2(_06634_),
    .B1(_06636_),
    .C1(_06446_),
    .X(_00390_));
 sky130_fd_sc_hd__clkbuf_4 _13906_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[0] ),
    .X(_06637_));
 sky130_fd_sc_hd__or2_1 _13907_ (.A(_06637_),
    .B(_05773_),
    .X(_06638_));
 sky130_fd_sc_hd__clkbuf_4 _13908_ (.A(_05260_),
    .X(_06639_));
 sky130_fd_sc_hd__o211a_1 _13909_ (.A1(_06618_),
    .A2(_06204_),
    .B1(_06638_),
    .C1(_06639_),
    .X(_00391_));
 sky130_fd_sc_hd__clkbuf_4 _13910_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[1] ),
    .X(_06640_));
 sky130_fd_sc_hd__buf_2 _13911_ (.A(_05772_),
    .X(_06641_));
 sky130_fd_sc_hd__or2_1 _13912_ (.A(_06640_),
    .B(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__o211a_1 _13913_ (.A1(_06622_),
    .A2(_06204_),
    .B1(_06642_),
    .C1(_06639_),
    .X(_00392_));
 sky130_fd_sc_hd__clkbuf_4 _13914_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[2] ),
    .X(_06643_));
 sky130_fd_sc_hd__or2_1 _13915_ (.A(_06643_),
    .B(_06641_),
    .X(_06644_));
 sky130_fd_sc_hd__o211a_1 _13916_ (.A1(_06624_),
    .A2(_06204_),
    .B1(_06644_),
    .C1(_06639_),
    .X(_00393_));
 sky130_fd_sc_hd__clkbuf_4 _13917_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[3] ),
    .X(_06645_));
 sky130_fd_sc_hd__or2_1 _13918_ (.A(_06645_),
    .B(_06641_),
    .X(_06646_));
 sky130_fd_sc_hd__o211a_1 _13919_ (.A1(_06626_),
    .A2(_06204_),
    .B1(_06646_),
    .C1(_06639_),
    .X(_00394_));
 sky130_fd_sc_hd__clkbuf_4 _13920_ (.A(_05755_),
    .X(_06647_));
 sky130_fd_sc_hd__clkbuf_4 _13921_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[4] ),
    .X(_06648_));
 sky130_fd_sc_hd__or2_1 _13922_ (.A(_06648_),
    .B(_06641_),
    .X(_06649_));
 sky130_fd_sc_hd__o211a_1 _13923_ (.A1(_06628_),
    .A2(_06647_),
    .B1(_06649_),
    .C1(_06639_),
    .X(_00395_));
 sky130_fd_sc_hd__clkbuf_4 _13924_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[5] ),
    .X(_06650_));
 sky130_fd_sc_hd__or2_1 _13925_ (.A(_06650_),
    .B(_06641_),
    .X(_06651_));
 sky130_fd_sc_hd__o211a_1 _13926_ (.A1(_06630_),
    .A2(_06647_),
    .B1(_06651_),
    .C1(_06639_),
    .X(_00396_));
 sky130_fd_sc_hd__clkbuf_4 _13927_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[6] ),
    .X(_06652_));
 sky130_fd_sc_hd__or2_1 _13928_ (.A(_06652_),
    .B(_06641_),
    .X(_06653_));
 sky130_fd_sc_hd__o211a_1 _13929_ (.A1(_06632_),
    .A2(_06647_),
    .B1(_06653_),
    .C1(_06639_),
    .X(_00397_));
 sky130_fd_sc_hd__or2_1 _13930_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[7] ),
    .B(_06641_),
    .X(_06654_));
 sky130_fd_sc_hd__o211a_1 _13931_ (.A1(_06635_),
    .A2(_06647_),
    .B1(_06654_),
    .C1(_06639_),
    .X(_00398_));
 sky130_fd_sc_hd__a21o_1 _13932_ (.A1(_06637_),
    .A2(_06618_),
    .B1(_05328_),
    .X(_06655_));
 sky130_fd_sc_hd__o211a_1 _13933_ (.A1(net1078),
    .A2(_05788_),
    .B1(_06655_),
    .C1(_06639_),
    .X(_00399_));
 sky130_fd_sc_hd__and4_1 _13934_ (.A(_06640_),
    .B(_06622_),
    .C(_06637_),
    .D(_06618_),
    .X(_06656_));
 sky130_fd_sc_hd__a22o_1 _13935_ (.A1(_06622_),
    .A2(_06637_),
    .B1(_06618_),
    .B2(_06640_),
    .X(_06657_));
 sky130_fd_sc_hd__or3b_1 _13936_ (.A(_05406_),
    .B(_06656_),
    .C_N(_06657_),
    .X(_06658_));
 sky130_fd_sc_hd__nand2_1 _13937_ (.A(net1000),
    .B(_05403_),
    .Y(_06659_));
 sky130_fd_sc_hd__a21oi_1 _13938_ (.A1(_06658_),
    .A2(_06659_),
    .B1(_05440_),
    .Y(_00400_));
 sky130_fd_sc_hd__buf_4 _13939_ (.A(_05787_),
    .X(_06660_));
 sky130_fd_sc_hd__nand4_2 _13940_ (.A(_06624_),
    .B(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[1] ),
    .C(_06622_),
    .D(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[0] ),
    .Y(_06661_));
 sky130_fd_sc_hd__or2_1 _13941_ (.A(_06656_),
    .B(_06661_),
    .X(_06662_));
 sky130_fd_sc_hd__a22o_1 _13942_ (.A1(_06640_),
    .A2(_06622_),
    .B1(_06637_),
    .B2(_06624_),
    .X(_06663_));
 sky130_fd_sc_hd__nand2_1 _13943_ (.A(_06656_),
    .B(_06661_),
    .Y(_06664_));
 sky130_fd_sc_hd__and2_1 _13944_ (.A(_06643_),
    .B(_06618_),
    .X(_06665_));
 sky130_fd_sc_hd__a31o_1 _13945_ (.A1(_06662_),
    .A2(_06663_),
    .A3(_06664_),
    .B1(_06665_),
    .X(_06666_));
 sky130_fd_sc_hd__nand4_2 _13946_ (.A(_06662_),
    .B(_06663_),
    .C(_06664_),
    .D(_06665_),
    .Y(_06667_));
 sky130_fd_sc_hd__a21o_1 _13947_ (.A1(_06666_),
    .A2(_06667_),
    .B1(_05328_),
    .X(_06668_));
 sky130_fd_sc_hd__o211a_1 _13948_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[2] ),
    .A2(_06660_),
    .B1(_06668_),
    .C1(_06639_),
    .X(_00401_));
 sky130_fd_sc_hd__a22oi_1 _13949_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[2] ),
    .A2(_06622_),
    .B1(_06618_),
    .B2(_06645_),
    .Y(_06669_));
 sky130_fd_sc_hd__and4_1 _13950_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[3] ),
    .B(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[2] ),
    .C(_06622_),
    .D(\top_inst.grid_inst.data_path_wires[3][0] ),
    .X(_06670_));
 sky130_fd_sc_hd__nor2_1 _13951_ (.A(_06669_),
    .B(_06670_),
    .Y(_06671_));
 sky130_fd_sc_hd__and4_1 _13952_ (.A(\top_inst.grid_inst.data_path_wires[3][3] ),
    .B(\top_inst.grid_inst.data_path_wires[3][2] ),
    .C(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[0] ),
    .X(_06672_));
 sky130_fd_sc_hd__nand2_1 _13953_ (.A(_06661_),
    .B(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__a22o_1 _13954_ (.A1(_06624_),
    .A2(_06640_),
    .B1(_06637_),
    .B2(_06626_),
    .X(_06674_));
 sky130_fd_sc_hd__or2_1 _13955_ (.A(_06661_),
    .B(_06672_),
    .X(_06675_));
 sky130_fd_sc_hd__and4_1 _13956_ (.A(_06671_),
    .B(_06673_),
    .C(_06674_),
    .D(_06675_),
    .X(_06676_));
 sky130_fd_sc_hd__a31o_1 _13957_ (.A1(_06673_),
    .A2(_06674_),
    .A3(_06675_),
    .B1(_06671_),
    .X(_06677_));
 sky130_fd_sc_hd__or2b_1 _13958_ (.A(_06676_),
    .B_N(_06677_),
    .X(_06678_));
 sky130_fd_sc_hd__xnor2_1 _13959_ (.A(_06667_),
    .B(_06678_),
    .Y(_06679_));
 sky130_fd_sc_hd__nand2_1 _13960_ (.A(_06664_),
    .B(_06679_),
    .Y(_06680_));
 sky130_fd_sc_hd__or2_1 _13961_ (.A(_06664_),
    .B(_06679_),
    .X(_06681_));
 sky130_fd_sc_hd__buf_6 _13962_ (.A(_05327_),
    .X(_06682_));
 sky130_fd_sc_hd__a21o_1 _13963_ (.A1(_06680_),
    .A2(_06681_),
    .B1(_06682_),
    .X(_06683_));
 sky130_fd_sc_hd__clkbuf_4 _13964_ (.A(_05260_),
    .X(_06684_));
 sky130_fd_sc_hd__o211a_1 _13965_ (.A1(net1072),
    .A2(_06660_),
    .B1(_06683_),
    .C1(_06684_),
    .X(_00402_));
 sky130_fd_sc_hd__inv_2 _13966_ (.A(_06672_),
    .Y(_06685_));
 sky130_fd_sc_hd__nand4_1 _13967_ (.A(\top_inst.grid_inst.data_path_wires[3][4] ),
    .B(\top_inst.grid_inst.data_path_wires[3][3] ),
    .C(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[0] ),
    .Y(_06686_));
 sky130_fd_sc_hd__a22o_1 _13968_ (.A1(\top_inst.grid_inst.data_path_wires[3][3] ),
    .A2(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[3][4] ),
    .X(_06687_));
 sky130_fd_sc_hd__nand2_1 _13969_ (.A(_06686_),
    .B(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__xor2_1 _13970_ (.A(_06670_),
    .B(_06688_),
    .X(_06689_));
 sky130_fd_sc_hd__xnor2_1 _13971_ (.A(_06685_),
    .B(_06689_),
    .Y(_06690_));
 sky130_fd_sc_hd__nand2_1 _13972_ (.A(_06643_),
    .B(_06624_),
    .Y(_06691_));
 sky130_fd_sc_hd__and3_1 _13973_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[3] ),
    .C(\top_inst.grid_inst.data_path_wires[3][1] ),
    .X(_06692_));
 sky130_fd_sc_hd__a22o_1 _13974_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[3] ),
    .A2(\top_inst.grid_inst.data_path_wires[3][1] ),
    .B1(\top_inst.grid_inst.data_path_wires[3][0] ),
    .B2(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[4] ),
    .X(_06693_));
 sky130_fd_sc_hd__a21bo_1 _13975_ (.A1(_06618_),
    .A2(_06692_),
    .B1_N(_06693_),
    .X(_06694_));
 sky130_fd_sc_hd__xor2_1 _13976_ (.A(_06691_),
    .B(_06694_),
    .X(_06695_));
 sky130_fd_sc_hd__xnor2_1 _13977_ (.A(_06690_),
    .B(_06695_),
    .Y(_06696_));
 sky130_fd_sc_hd__xnor2_1 _13978_ (.A(_06676_),
    .B(_06696_),
    .Y(_06697_));
 sky130_fd_sc_hd__xnor2_1 _13979_ (.A(_06675_),
    .B(_06697_),
    .Y(_06698_));
 sky130_fd_sc_hd__o21ai_1 _13980_ (.A1(_06667_),
    .A2(_06678_),
    .B1(_06681_),
    .Y(_06699_));
 sky130_fd_sc_hd__xnor2_1 _13981_ (.A(_06698_),
    .B(_06699_),
    .Y(_06700_));
 sky130_fd_sc_hd__buf_8 _13982_ (.A(_05311_),
    .X(_06701_));
 sky130_fd_sc_hd__mux2_1 _13983_ (.A0(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[4] ),
    .A1(_06700_),
    .S(_06701_),
    .X(_06702_));
 sky130_fd_sc_hd__and2_1 _13984_ (.A(_06364_),
    .B(_06702_),
    .X(_06703_));
 sky130_fd_sc_hd__clkbuf_1 _13985_ (.A(_06703_),
    .X(_00403_));
 sky130_fd_sc_hd__or2b_1 _13986_ (.A(_06698_),
    .B_N(_06699_),
    .X(_06704_));
 sky130_fd_sc_hd__nand2_1 _13987_ (.A(_06676_),
    .B(_06696_),
    .Y(_06705_));
 sky130_fd_sc_hd__or2_1 _13988_ (.A(_06675_),
    .B(_06697_),
    .X(_06706_));
 sky130_fd_sc_hd__or2b_1 _13989_ (.A(_06690_),
    .B_N(_06695_),
    .X(_06707_));
 sky130_fd_sc_hd__nand2_1 _13990_ (.A(_06650_),
    .B(_06618_),
    .Y(_06708_));
 sky130_fd_sc_hd__a22o_1 _13991_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[3] ),
    .A2(\top_inst.grid_inst.data_path_wires[3][2] ),
    .B1(\top_inst.grid_inst.data_path_wires[3][1] ),
    .B2(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[4] ),
    .X(_06709_));
 sky130_fd_sc_hd__nand4_1 _13992_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[3] ),
    .C(\top_inst.grid_inst.data_path_wires[3][2] ),
    .D(\top_inst.grid_inst.data_path_wires[3][1] ),
    .Y(_06710_));
 sky130_fd_sc_hd__a22oi_2 _13993_ (.A1(_06626_),
    .A2(_06643_),
    .B1(_06709_),
    .B2(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__and4_1 _13994_ (.A(_06626_),
    .B(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[2] ),
    .C(_06709_),
    .D(_06710_),
    .X(_06712_));
 sky130_fd_sc_hd__nor2_1 _13995_ (.A(_06711_),
    .B(_06712_),
    .Y(_06713_));
 sky130_fd_sc_hd__xnor2_2 _13996_ (.A(_06708_),
    .B(_06713_),
    .Y(_06714_));
 sky130_fd_sc_hd__and4_1 _13997_ (.A(_06628_),
    .B(_06626_),
    .C(_06640_),
    .D(_06637_),
    .X(_06715_));
 sky130_fd_sc_hd__a32o_1 _13998_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[2] ),
    .A2(_06624_),
    .A3(_06693_),
    .B1(_06692_),
    .B2(\top_inst.grid_inst.data_path_wires[3][0] ),
    .X(_06716_));
 sky130_fd_sc_hd__and4_1 _13999_ (.A(\top_inst.grid_inst.data_path_wires[3][5] ),
    .B(\top_inst.grid_inst.data_path_wires[3][4] ),
    .C(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[0] ),
    .X(_06717_));
 sky130_fd_sc_hd__a22oi_1 _14000_ (.A1(\top_inst.grid_inst.data_path_wires[3][4] ),
    .A2(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[3][5] ),
    .Y(_06718_));
 sky130_fd_sc_hd__nor2_1 _14001_ (.A(_06717_),
    .B(_06718_),
    .Y(_06719_));
 sky130_fd_sc_hd__xor2_1 _14002_ (.A(_06716_),
    .B(_06719_),
    .X(_06720_));
 sky130_fd_sc_hd__xnor2_1 _14003_ (.A(_06715_),
    .B(_06720_),
    .Y(_06721_));
 sky130_fd_sc_hd__xor2_1 _14004_ (.A(_06714_),
    .B(_06721_),
    .X(_06722_));
 sky130_fd_sc_hd__xor2_1 _14005_ (.A(_06707_),
    .B(_06722_),
    .X(_06723_));
 sky130_fd_sc_hd__nor2_1 _14006_ (.A(_06685_),
    .B(_06689_),
    .Y(_06724_));
 sky130_fd_sc_hd__a31o_1 _14007_ (.A1(_06670_),
    .A2(_06686_),
    .A3(_06687_),
    .B1(_06724_),
    .X(_06725_));
 sky130_fd_sc_hd__xnor2_1 _14008_ (.A(_06723_),
    .B(_06725_),
    .Y(_06726_));
 sky130_fd_sc_hd__a21oi_1 _14009_ (.A1(_06705_),
    .A2(_06706_),
    .B1(_06726_),
    .Y(_06727_));
 sky130_fd_sc_hd__and3_1 _14010_ (.A(_06705_),
    .B(_06706_),
    .C(_06726_),
    .X(_06728_));
 sky130_fd_sc_hd__or2_1 _14011_ (.A(_06727_),
    .B(_06728_),
    .X(_06729_));
 sky130_fd_sc_hd__or2_1 _14012_ (.A(_06704_),
    .B(_06729_),
    .X(_06730_));
 sky130_fd_sc_hd__a21oi_1 _14013_ (.A1(_06704_),
    .A2(_06729_),
    .B1(_05399_),
    .Y(_06731_));
 sky130_fd_sc_hd__a22o_1 _14014_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[5] ),
    .A2(_06242_),
    .B1(_06730_),
    .B2(_06731_),
    .X(_06732_));
 sky130_fd_sc_hd__and2_1 _14015_ (.A(_06364_),
    .B(_06732_),
    .X(_06733_));
 sky130_fd_sc_hd__clkbuf_1 _14016_ (.A(_06733_),
    .X(_00404_));
 sky130_fd_sc_hd__buf_8 _14017_ (.A(_05633_),
    .X(_06734_));
 sky130_fd_sc_hd__nand2_1 _14018_ (.A(_06716_),
    .B(_06719_),
    .Y(_06735_));
 sky130_fd_sc_hd__nand2_1 _14019_ (.A(_06715_),
    .B(_06720_),
    .Y(_06736_));
 sky130_fd_sc_hd__inv_2 _14020_ (.A(_06714_),
    .Y(_06737_));
 sky130_fd_sc_hd__nor2_1 _14021_ (.A(_06737_),
    .B(_06721_),
    .Y(_06738_));
 sky130_fd_sc_hd__or3_2 _14022_ (.A(_06708_),
    .B(_06711_),
    .C(_06712_),
    .X(_06739_));
 sky130_fd_sc_hd__a22o_1 _14023_ (.A1(_06650_),
    .A2(_06622_),
    .B1(_06618_),
    .B2(_06652_),
    .X(_06740_));
 sky130_fd_sc_hd__nand4_4 _14024_ (.A(_06652_),
    .B(_06650_),
    .C(_06622_),
    .D(\top_inst.grid_inst.data_path_wires[3][0] ),
    .Y(_06741_));
 sky130_fd_sc_hd__nand2_1 _14025_ (.A(_06740_),
    .B(_06741_),
    .Y(_06742_));
 sky130_fd_sc_hd__a22o_1 _14026_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[3] ),
    .A2(\top_inst.grid_inst.data_path_wires[3][3] ),
    .B1(\top_inst.grid_inst.data_path_wires[3][2] ),
    .B2(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[4] ),
    .X(_06743_));
 sky130_fd_sc_hd__nand4_2 _14027_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[3] ),
    .C(\top_inst.grid_inst.data_path_wires[3][3] ),
    .D(_06624_),
    .Y(_06744_));
 sky130_fd_sc_hd__a22o_1 _14028_ (.A1(_06628_),
    .A2(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[2] ),
    .B1(_06743_),
    .B2(_06744_),
    .X(_06745_));
 sky130_fd_sc_hd__nand4_1 _14029_ (.A(_06628_),
    .B(_06643_),
    .C(_06743_),
    .D(_06744_),
    .Y(_06746_));
 sky130_fd_sc_hd__nand2_1 _14030_ (.A(_06745_),
    .B(_06746_),
    .Y(_06747_));
 sky130_fd_sc_hd__xnor2_2 _14031_ (.A(_06742_),
    .B(_06747_),
    .Y(_06748_));
 sky130_fd_sc_hd__xnor2_2 _14032_ (.A(_06739_),
    .B(_06748_),
    .Y(_06749_));
 sky130_fd_sc_hd__a21o_1 _14033_ (.A1(_06624_),
    .A2(_06692_),
    .B1(_06712_),
    .X(_06750_));
 sky130_fd_sc_hd__and4_2 _14034_ (.A(\top_inst.grid_inst.data_path_wires[3][6] ),
    .B(\top_inst.grid_inst.data_path_wires[3][5] ),
    .C(_06640_),
    .D(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[0] ),
    .X(_06751_));
 sky130_fd_sc_hd__a22oi_1 _14035_ (.A1(_06630_),
    .A2(_06640_),
    .B1(_06637_),
    .B2(\top_inst.grid_inst.data_path_wires[3][6] ),
    .Y(_06752_));
 sky130_fd_sc_hd__nor2_1 _14036_ (.A(_06751_),
    .B(_06752_),
    .Y(_06753_));
 sky130_fd_sc_hd__xor2_2 _14037_ (.A(_06750_),
    .B(_06753_),
    .X(_06754_));
 sky130_fd_sc_hd__xnor2_2 _14038_ (.A(_06717_),
    .B(_06754_),
    .Y(_06755_));
 sky130_fd_sc_hd__xnor2_2 _14039_ (.A(_06749_),
    .B(_06755_),
    .Y(_06756_));
 sky130_fd_sc_hd__xor2_1 _14040_ (.A(_06738_),
    .B(_06756_),
    .X(_06757_));
 sky130_fd_sc_hd__a21oi_2 _14041_ (.A1(_06735_),
    .A2(_06736_),
    .B1(_06757_),
    .Y(_06758_));
 sky130_fd_sc_hd__and3_1 _14042_ (.A(_06735_),
    .B(_06736_),
    .C(_06757_),
    .X(_06759_));
 sky130_fd_sc_hd__nor2_1 _14043_ (.A(_06707_),
    .B(_06722_),
    .Y(_06760_));
 sky130_fd_sc_hd__a21oi_1 _14044_ (.A1(_06723_),
    .A2(_06725_),
    .B1(_06760_),
    .Y(_06761_));
 sky130_fd_sc_hd__nor3_1 _14045_ (.A(_06758_),
    .B(_06759_),
    .C(_06761_),
    .Y(_06762_));
 sky130_fd_sc_hd__o21a_1 _14046_ (.A1(_06758_),
    .A2(_06759_),
    .B1(_06761_),
    .X(_06763_));
 sky130_fd_sc_hd__o21ba_1 _14047_ (.A1(_06704_),
    .A2(_06728_),
    .B1_N(_06727_),
    .X(_06764_));
 sky130_fd_sc_hd__nor3_1 _14048_ (.A(_06762_),
    .B(_06763_),
    .C(_06764_),
    .Y(_06765_));
 sky130_fd_sc_hd__o21a_1 _14049_ (.A1(_06762_),
    .A2(_06763_),
    .B1(_06764_),
    .X(_06766_));
 sky130_fd_sc_hd__nand2_1 _14050_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[6] ),
    .B(_05406_),
    .Y(_06767_));
 sky130_fd_sc_hd__o31a_1 _14051_ (.A1(_06734_),
    .A2(_06765_),
    .A3(_06766_),
    .B1(_06767_),
    .X(_06768_));
 sky130_fd_sc_hd__nor2_1 _14052_ (.A(_05632_),
    .B(_06768_),
    .Y(_00405_));
 sky130_fd_sc_hd__nor2_1 _14053_ (.A(_06742_),
    .B(_06747_),
    .Y(_06769_));
 sky130_fd_sc_hd__nand2_1 _14054_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[6] ),
    .B(\top_inst.grid_inst.data_path_wires[3][1] ),
    .Y(_06770_));
 sky130_fd_sc_hd__or2b_1 _14055_ (.A(\top_inst.grid_inst.data_path_wires[3][0] ),
    .B_N(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[7] ),
    .X(_06771_));
 sky130_fd_sc_hd__xnor2_2 _14056_ (.A(_06770_),
    .B(_06771_),
    .Y(_06772_));
 sky130_fd_sc_hd__nand2_1 _14057_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[5] ),
    .B(_06624_),
    .Y(_06773_));
 sky130_fd_sc_hd__xnor2_2 _14058_ (.A(_06772_),
    .B(_06773_),
    .Y(_06774_));
 sky130_fd_sc_hd__xor2_2 _14059_ (.A(_06741_),
    .B(_06774_),
    .X(_06775_));
 sky130_fd_sc_hd__a22o_1 _14060_ (.A1(\top_inst.grid_inst.data_path_wires[3][4] ),
    .A2(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[3] ),
    .B1(_06626_),
    .B2(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[4] ),
    .X(_06776_));
 sky130_fd_sc_hd__nand4_4 _14061_ (.A(_06648_),
    .B(_06628_),
    .C(_06645_),
    .D(_06626_),
    .Y(_06777_));
 sky130_fd_sc_hd__a22o_1 _14062_ (.A1(_06630_),
    .A2(_06643_),
    .B1(_06776_),
    .B2(_06777_),
    .X(_06778_));
 sky130_fd_sc_hd__nand4_2 _14063_ (.A(_06630_),
    .B(_06643_),
    .C(_06776_),
    .D(_06777_),
    .Y(_06779_));
 sky130_fd_sc_hd__nand2_1 _14064_ (.A(_06778_),
    .B(_06779_),
    .Y(_06780_));
 sky130_fd_sc_hd__xnor2_2 _14065_ (.A(_06775_),
    .B(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__xnor2_2 _14066_ (.A(_06769_),
    .B(_06781_),
    .Y(_06782_));
 sky130_fd_sc_hd__nand2_1 _14067_ (.A(_06744_),
    .B(_06746_),
    .Y(_06783_));
 sky130_fd_sc_hd__a22o_1 _14068_ (.A1(\top_inst.grid_inst.data_path_wires[3][6] ),
    .A2(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[3][7] ),
    .X(_06784_));
 sky130_fd_sc_hd__and3_1 _14069_ (.A(\top_inst.grid_inst.data_path_wires[3][7] ),
    .B(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[1] ),
    .C(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[0] ),
    .X(_06785_));
 sky130_fd_sc_hd__nand2_1 _14070_ (.A(\top_inst.grid_inst.data_path_wires[3][6] ),
    .B(_06785_),
    .Y(_06786_));
 sky130_fd_sc_hd__and3_1 _14071_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[7] ),
    .B(_06784_),
    .C(_06786_),
    .X(_06787_));
 sky130_fd_sc_hd__a21oi_1 _14072_ (.A1(_06784_),
    .A2(_06786_),
    .B1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[7] ),
    .Y(_06788_));
 sky130_fd_sc_hd__or2_1 _14073_ (.A(_06787_),
    .B(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__xnor2_2 _14074_ (.A(_06783_),
    .B(_06789_),
    .Y(_06790_));
 sky130_fd_sc_hd__xnor2_2 _14075_ (.A(_06751_),
    .B(_06790_),
    .Y(_06791_));
 sky130_fd_sc_hd__xor2_2 _14076_ (.A(_06782_),
    .B(_06791_),
    .X(_06792_));
 sky130_fd_sc_hd__or2_1 _14077_ (.A(_06739_),
    .B(_06748_),
    .X(_06793_));
 sky130_fd_sc_hd__o21ai_2 _14078_ (.A1(_06749_),
    .A2(_06755_),
    .B1(_06793_),
    .Y(_06794_));
 sky130_fd_sc_hd__xnor2_2 _14079_ (.A(_06792_),
    .B(_06794_),
    .Y(_06795_));
 sky130_fd_sc_hd__and2_1 _14080_ (.A(_06750_),
    .B(_06753_),
    .X(_06796_));
 sky130_fd_sc_hd__a21o_1 _14081_ (.A1(_06717_),
    .A2(_06754_),
    .B1(_06796_),
    .X(_06797_));
 sky130_fd_sc_hd__xnor2_2 _14082_ (.A(_06795_),
    .B(_06797_),
    .Y(_06798_));
 sky130_fd_sc_hd__inv_2 _14083_ (.A(_06756_),
    .Y(_06799_));
 sky130_fd_sc_hd__a21oi_2 _14084_ (.A1(_06738_),
    .A2(_06799_),
    .B1(_06758_),
    .Y(_06800_));
 sky130_fd_sc_hd__xnor2_2 _14085_ (.A(_06798_),
    .B(_06800_),
    .Y(_06801_));
 sky130_fd_sc_hd__o21bai_2 _14086_ (.A1(_06763_),
    .A2(_06764_),
    .B1_N(_06762_),
    .Y(_06802_));
 sky130_fd_sc_hd__nor2_1 _14087_ (.A(_06801_),
    .B(_06802_),
    .Y(_06803_));
 sky130_fd_sc_hd__a21o_1 _14088_ (.A1(_06801_),
    .A2(_06802_),
    .B1(_05633_),
    .X(_06804_));
 sky130_fd_sc_hd__o2bb2a_1 _14089_ (.A1_N(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[7] ),
    .A2_N(_05634_),
    .B1(_06803_),
    .B2(_06804_),
    .X(_06805_));
 sky130_fd_sc_hd__nor2_1 _14090_ (.A(_05632_),
    .B(_06805_),
    .Y(_00406_));
 sky130_fd_sc_hd__and2b_1 _14091_ (.A_N(\top_inst.grid_inst.data_path_wires[3][1] ),
    .B(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[7] ),
    .X(_06806_));
 sky130_fd_sc_hd__a21oi_1 _14092_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[6] ),
    .A2(\top_inst.grid_inst.data_path_wires[3][2] ),
    .B1(_06806_),
    .Y(_06807_));
 sky130_fd_sc_hd__and3_1 _14093_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[6] ),
    .B(\top_inst.grid_inst.data_path_wires[3][2] ),
    .C(_06806_),
    .X(_06808_));
 sky130_fd_sc_hd__nor2_1 _14094_ (.A(_06807_),
    .B(_06808_),
    .Y(_06809_));
 sky130_fd_sc_hd__nand2_1 _14095_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[5] ),
    .B(_06626_),
    .Y(_06810_));
 sky130_fd_sc_hd__xnor2_2 _14096_ (.A(_06809_),
    .B(_06810_),
    .Y(_06811_));
 sky130_fd_sc_hd__nor2_1 _14097_ (.A(_06772_),
    .B(_06773_),
    .Y(_06812_));
 sky130_fd_sc_hd__o21ba_1 _14098_ (.A1(_06770_),
    .A2(_06771_),
    .B1_N(_06812_),
    .X(_06813_));
 sky130_fd_sc_hd__xnor2_2 _14099_ (.A(_06811_),
    .B(_06813_),
    .Y(_06814_));
 sky130_fd_sc_hd__a22o_1 _14100_ (.A1(_06648_),
    .A2(\top_inst.grid_inst.data_path_wires[3][4] ),
    .B1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[3][5] ),
    .X(_06815_));
 sky130_fd_sc_hd__nand4_1 _14101_ (.A(\top_inst.grid_inst.data_path_wires[3][5] ),
    .B(_06648_),
    .C(_06628_),
    .D(_06645_),
    .Y(_06816_));
 sky130_fd_sc_hd__a22oi_1 _14102_ (.A1(_06632_),
    .A2(_06643_),
    .B1(_06815_),
    .B2(_06816_),
    .Y(_06817_));
 sky130_fd_sc_hd__and4_1 _14103_ (.A(_06632_),
    .B(_06643_),
    .C(_06815_),
    .D(_06816_),
    .X(_06818_));
 sky130_fd_sc_hd__or2_1 _14104_ (.A(_06817_),
    .B(_06818_),
    .X(_06819_));
 sky130_fd_sc_hd__xnor2_2 _14105_ (.A(_06814_),
    .B(_06819_),
    .Y(_06820_));
 sky130_fd_sc_hd__and3_1 _14106_ (.A(_06775_),
    .B(_06778_),
    .C(_06779_),
    .X(_06821_));
 sky130_fd_sc_hd__o21ba_1 _14107_ (.A1(_06741_),
    .A2(_06774_),
    .B1_N(_06821_),
    .X(_06822_));
 sky130_fd_sc_hd__xnor2_2 _14108_ (.A(_06820_),
    .B(_06822_),
    .Y(_06823_));
 sky130_fd_sc_hd__and2_1 _14109_ (.A(_06632_),
    .B(_06785_),
    .X(_06824_));
 sky130_fd_sc_hd__o21ai_4 _14110_ (.A1(_06640_),
    .A2(_06637_),
    .B1(\top_inst.grid_inst.data_path_wires[3][7] ),
    .Y(_06825_));
 sky130_fd_sc_hd__or2_1 _14111_ (.A(_06785_),
    .B(_06825_),
    .X(_06826_));
 sky130_fd_sc_hd__a21o_1 _14112_ (.A1(_06777_),
    .A2(_06779_),
    .B1(_06826_),
    .X(_06827_));
 sky130_fd_sc_hd__nand3_1 _14113_ (.A(_06777_),
    .B(_06779_),
    .C(_06826_),
    .Y(_06828_));
 sky130_fd_sc_hd__o211a_1 _14114_ (.A1(_06824_),
    .A2(_06787_),
    .B1(_06827_),
    .C1(_06828_),
    .X(_06829_));
 sky130_fd_sc_hd__nor2_1 _14115_ (.A(_06824_),
    .B(_06787_),
    .Y(_06830_));
 sky130_fd_sc_hd__a21boi_1 _14116_ (.A1(_06827_),
    .A2(_06828_),
    .B1_N(_06830_),
    .Y(_06831_));
 sky130_fd_sc_hd__nor2_1 _14117_ (.A(_06829_),
    .B(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__xnor2_2 _14118_ (.A(_06823_),
    .B(_06832_),
    .Y(_06833_));
 sky130_fd_sc_hd__nand2_1 _14119_ (.A(_06769_),
    .B(_06781_),
    .Y(_06834_));
 sky130_fd_sc_hd__o21a_1 _14120_ (.A1(_06782_),
    .A2(_06791_),
    .B1(_06834_),
    .X(_06835_));
 sky130_fd_sc_hd__xnor2_2 _14121_ (.A(_06833_),
    .B(_06835_),
    .Y(_06836_));
 sky130_fd_sc_hd__or2b_1 _14122_ (.A(_06789_),
    .B_N(_06783_),
    .X(_06837_));
 sky130_fd_sc_hd__a21boi_2 _14123_ (.A1(_06751_),
    .A2(_06790_),
    .B1_N(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__xnor2_2 _14124_ (.A(_06836_),
    .B(_06838_),
    .Y(_06839_));
 sky130_fd_sc_hd__or2b_1 _14125_ (.A(_06795_),
    .B_N(_06797_),
    .X(_06840_));
 sky130_fd_sc_hd__a21boi_2 _14126_ (.A1(_06792_),
    .A2(_06794_),
    .B1_N(_06840_),
    .Y(_06841_));
 sky130_fd_sc_hd__xnor2_2 _14127_ (.A(_06839_),
    .B(_06841_),
    .Y(_06842_));
 sky130_fd_sc_hd__or2b_1 _14128_ (.A(_06800_),
    .B_N(_06798_),
    .X(_06843_));
 sky130_fd_sc_hd__a21boi_2 _14129_ (.A1(_06801_),
    .A2(_06802_),
    .B1_N(_06843_),
    .Y(_06844_));
 sky130_fd_sc_hd__nor2_1 _14130_ (.A(_06842_),
    .B(_06844_),
    .Y(_06845_));
 sky130_fd_sc_hd__a21o_1 _14131_ (.A1(_06842_),
    .A2(_06844_),
    .B1(_05633_),
    .X(_06846_));
 sky130_fd_sc_hd__o2bb2a_1 _14132_ (.A1_N(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[8] ),
    .A2_N(_05634_),
    .B1(_06845_),
    .B2(_06846_),
    .X(_06847_));
 sky130_fd_sc_hd__nor2_1 _14133_ (.A(_05632_),
    .B(_06847_),
    .Y(_00407_));
 sky130_fd_sc_hd__buf_4 _14134_ (.A(_05732_),
    .X(_06848_));
 sky130_fd_sc_hd__and2b_1 _14135_ (.A_N(\top_inst.grid_inst.data_path_wires[3][2] ),
    .B(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[7] ),
    .X(_06849_));
 sky130_fd_sc_hd__a21oi_1 _14136_ (.A1(_06652_),
    .A2(_06626_),
    .B1(_06849_),
    .Y(_06850_));
 sky130_fd_sc_hd__and3_1 _14137_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[6] ),
    .B(\top_inst.grid_inst.data_path_wires[3][3] ),
    .C(_06849_),
    .X(_06851_));
 sky130_fd_sc_hd__nor2_1 _14138_ (.A(_06850_),
    .B(_06851_),
    .Y(_06852_));
 sky130_fd_sc_hd__nand2_1 _14139_ (.A(_06650_),
    .B(_06628_),
    .Y(_06853_));
 sky130_fd_sc_hd__xnor2_1 _14140_ (.A(_06852_),
    .B(_06853_),
    .Y(_06854_));
 sky130_fd_sc_hd__o21ba_1 _14141_ (.A1(_06807_),
    .A2(_06810_),
    .B1_N(_06808_),
    .X(_06855_));
 sky130_fd_sc_hd__xor2_1 _14142_ (.A(_06854_),
    .B(_06855_),
    .X(_06856_));
 sky130_fd_sc_hd__a22oi_2 _14143_ (.A1(_06630_),
    .A2(_06648_),
    .B1(_06645_),
    .B2(_06632_),
    .Y(_06857_));
 sky130_fd_sc_hd__and4_1 _14144_ (.A(\top_inst.grid_inst.data_path_wires[3][6] ),
    .B(\top_inst.grid_inst.data_path_wires[3][5] ),
    .C(_06648_),
    .D(_06645_),
    .X(_06858_));
 sky130_fd_sc_hd__nor2_1 _14145_ (.A(_06857_),
    .B(_06858_),
    .Y(_06859_));
 sky130_fd_sc_hd__nand2_2 _14146_ (.A(_06635_),
    .B(_06643_),
    .Y(_06860_));
 sky130_fd_sc_hd__xor2_1 _14147_ (.A(_06859_),
    .B(_06860_),
    .X(_06861_));
 sky130_fd_sc_hd__xor2_1 _14148_ (.A(_06856_),
    .B(_06861_),
    .X(_06862_));
 sky130_fd_sc_hd__inv_2 _14149_ (.A(_06813_),
    .Y(_06863_));
 sky130_fd_sc_hd__or3b_1 _14150_ (.A(_06817_),
    .B(_06818_),
    .C_N(_06814_),
    .X(_06864_));
 sky130_fd_sc_hd__a21boi_1 _14151_ (.A1(_06811_),
    .A2(_06863_),
    .B1_N(_06864_),
    .Y(_06865_));
 sky130_fd_sc_hd__xnor2_1 _14152_ (.A(_06862_),
    .B(_06865_),
    .Y(_06866_));
 sky130_fd_sc_hd__and4_1 _14153_ (.A(_06630_),
    .B(_06648_),
    .C(_06628_),
    .D(_06645_),
    .X(_06867_));
 sky130_fd_sc_hd__nor2_1 _14154_ (.A(_06867_),
    .B(_06818_),
    .Y(_06868_));
 sky130_fd_sc_hd__nor2_1 _14155_ (.A(_06825_),
    .B(_06868_),
    .Y(_06869_));
 sky130_fd_sc_hd__and2_1 _14156_ (.A(_06825_),
    .B(_06868_),
    .X(_06870_));
 sky130_fd_sc_hd__nor2_1 _14157_ (.A(_06869_),
    .B(_06870_),
    .Y(_06871_));
 sky130_fd_sc_hd__xnor2_1 _14158_ (.A(_06866_),
    .B(_06871_),
    .Y(_06872_));
 sky130_fd_sc_hd__and2b_1 _14159_ (.A_N(_06822_),
    .B(_06820_),
    .X(_06873_));
 sky130_fd_sc_hd__a21oi_1 _14160_ (.A1(_06823_),
    .A2(_06832_),
    .B1(_06873_),
    .Y(_06874_));
 sky130_fd_sc_hd__xnor2_1 _14161_ (.A(_06872_),
    .B(_06874_),
    .Y(_06875_));
 sky130_fd_sc_hd__and3_1 _14162_ (.A(_06777_),
    .B(_06779_),
    .C(_06826_),
    .X(_06876_));
 sky130_fd_sc_hd__o21a_1 _14163_ (.A1(_06830_),
    .A2(_06876_),
    .B1(_06827_),
    .X(_06877_));
 sky130_fd_sc_hd__xnor2_1 _14164_ (.A(_06875_),
    .B(_06877_),
    .Y(_06878_));
 sky130_fd_sc_hd__or2_1 _14165_ (.A(_06833_),
    .B(_06835_),
    .X(_06879_));
 sky130_fd_sc_hd__o21a_1 _14166_ (.A1(_06836_),
    .A2(_06838_),
    .B1(_06879_),
    .X(_06880_));
 sky130_fd_sc_hd__nor2_1 _14167_ (.A(_06878_),
    .B(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__nand2_1 _14168_ (.A(_06878_),
    .B(_06880_),
    .Y(_06882_));
 sky130_fd_sc_hd__or2b_1 _14169_ (.A(_06881_),
    .B_N(_06882_),
    .X(_06883_));
 sky130_fd_sc_hd__nor2_1 _14170_ (.A(_06839_),
    .B(_06841_),
    .Y(_06884_));
 sky130_fd_sc_hd__o21bai_2 _14171_ (.A1(_06842_),
    .A2(_06844_),
    .B1_N(_06884_),
    .Y(_06885_));
 sky130_fd_sc_hd__xnor2_1 _14172_ (.A(_06883_),
    .B(_06885_),
    .Y(_06886_));
 sky130_fd_sc_hd__or2_1 _14173_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[9] ),
    .B(_06168_),
    .X(_06887_));
 sky130_fd_sc_hd__o211a_1 _14174_ (.A1(_06848_),
    .A2(_06886_),
    .B1(_06887_),
    .C1(_06684_),
    .X(_00408_));
 sky130_fd_sc_hd__or2b_1 _14175_ (.A(_06855_),
    .B_N(_06854_),
    .X(_06888_));
 sky130_fd_sc_hd__o21a_1 _14176_ (.A1(_06856_),
    .A2(_06861_),
    .B1(_06888_),
    .X(_06889_));
 sky130_fd_sc_hd__and2b_1 _14177_ (.A_N(\top_inst.grid_inst.data_path_wires[3][3] ),
    .B(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[7] ),
    .X(_06890_));
 sky130_fd_sc_hd__a21oi_1 _14178_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[6] ),
    .A2(_06628_),
    .B1(_06890_),
    .Y(_06891_));
 sky130_fd_sc_hd__and3_1 _14179_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[6] ),
    .B(\top_inst.grid_inst.data_path_wires[3][4] ),
    .C(_06890_),
    .X(_06892_));
 sky130_fd_sc_hd__nor2_1 _14180_ (.A(_06891_),
    .B(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__nand2_1 _14181_ (.A(_06650_),
    .B(_06630_),
    .Y(_06894_));
 sky130_fd_sc_hd__xnor2_1 _14182_ (.A(_06893_),
    .B(_06894_),
    .Y(_06895_));
 sky130_fd_sc_hd__o21ba_1 _14183_ (.A1(_06850_),
    .A2(_06853_),
    .B1_N(_06851_),
    .X(_06896_));
 sky130_fd_sc_hd__xor2_1 _14184_ (.A(_06895_),
    .B(_06896_),
    .X(_06897_));
 sky130_fd_sc_hd__and3_2 _14185_ (.A(\top_inst.grid_inst.data_path_wires[3][7] ),
    .B(_06648_),
    .C(_06645_),
    .X(_06898_));
 sky130_fd_sc_hd__a22oi_1 _14186_ (.A1(\top_inst.grid_inst.data_path_wires[3][6] ),
    .A2(_06648_),
    .B1(_06645_),
    .B2(_06635_),
    .Y(_06899_));
 sky130_fd_sc_hd__a21oi_1 _14187_ (.A1(_06632_),
    .A2(_06898_),
    .B1(_06899_),
    .Y(_06900_));
 sky130_fd_sc_hd__xnor2_1 _14188_ (.A(_06860_),
    .B(_06900_),
    .Y(_06901_));
 sky130_fd_sc_hd__xnor2_1 _14189_ (.A(_06897_),
    .B(_06901_),
    .Y(_06902_));
 sky130_fd_sc_hd__and2b_1 _14190_ (.A_N(_06889_),
    .B(_06902_),
    .X(_06903_));
 sky130_fd_sc_hd__and2b_1 _14191_ (.A_N(_06902_),
    .B(_06889_),
    .X(_06904_));
 sky130_fd_sc_hd__nor2_1 _14192_ (.A(_06903_),
    .B(_06904_),
    .Y(_06905_));
 sky130_fd_sc_hd__o21ba_1 _14193_ (.A1(_06857_),
    .A2(_06860_),
    .B1_N(_06858_),
    .X(_06906_));
 sky130_fd_sc_hd__nor2_1 _14194_ (.A(_06825_),
    .B(_06906_),
    .Y(_06907_));
 sky130_fd_sc_hd__and2_1 _14195_ (.A(_06825_),
    .B(_06906_),
    .X(_06908_));
 sky130_fd_sc_hd__nor2_1 _14196_ (.A(_06907_),
    .B(_06908_),
    .Y(_06909_));
 sky130_fd_sc_hd__xnor2_1 _14197_ (.A(_06905_),
    .B(_06909_),
    .Y(_06910_));
 sky130_fd_sc_hd__and2b_1 _14198_ (.A_N(_06865_),
    .B(_06862_),
    .X(_06911_));
 sky130_fd_sc_hd__a21oi_1 _14199_ (.A1(_06866_),
    .A2(_06871_),
    .B1(_06911_),
    .Y(_06912_));
 sky130_fd_sc_hd__xor2_1 _14200_ (.A(_06910_),
    .B(_06912_),
    .X(_06913_));
 sky130_fd_sc_hd__xnor2_1 _14201_ (.A(_06869_),
    .B(_06913_),
    .Y(_06914_));
 sky130_fd_sc_hd__or2_1 _14202_ (.A(_06872_),
    .B(_06874_),
    .X(_06915_));
 sky130_fd_sc_hd__o21a_1 _14203_ (.A1(_06875_),
    .A2(_06877_),
    .B1(_06915_),
    .X(_06916_));
 sky130_fd_sc_hd__nor2_1 _14204_ (.A(_06914_),
    .B(_06916_),
    .Y(_06917_));
 sky130_fd_sc_hd__and2_1 _14205_ (.A(_06914_),
    .B(_06916_),
    .X(_06918_));
 sky130_fd_sc_hd__or2_1 _14206_ (.A(_06917_),
    .B(_06918_),
    .X(_06919_));
 sky130_fd_sc_hd__a21oi_2 _14207_ (.A1(_06882_),
    .A2(_06885_),
    .B1(_06881_),
    .Y(_06920_));
 sky130_fd_sc_hd__nor2_1 _14208_ (.A(_06919_),
    .B(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__a21o_1 _14209_ (.A1(_06919_),
    .A2(_06920_),
    .B1(_06404_),
    .X(_06922_));
 sky130_fd_sc_hd__a2bb2o_1 _14210_ (.A1_N(_06921_),
    .A2_N(_06922_),
    .B1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[10] ),
    .B2(_05327_),
    .X(_06923_));
 sky130_fd_sc_hd__and2_1 _14211_ (.A(_06364_),
    .B(_06923_),
    .X(_06924_));
 sky130_fd_sc_hd__clkbuf_1 _14212_ (.A(_06924_),
    .X(_00409_));
 sky130_fd_sc_hd__and2b_1 _14213_ (.A_N(\top_inst.grid_inst.data_path_wires[3][4] ),
    .B(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[7] ),
    .X(_06925_));
 sky130_fd_sc_hd__a21oi_1 _14214_ (.A1(_06652_),
    .A2(\top_inst.grid_inst.data_path_wires[3][5] ),
    .B1(_06925_),
    .Y(_06926_));
 sky130_fd_sc_hd__and3_1 _14215_ (.A(_06652_),
    .B(\top_inst.grid_inst.data_path_wires[3][5] ),
    .C(_06925_),
    .X(_06927_));
 sky130_fd_sc_hd__nor2_1 _14216_ (.A(_06926_),
    .B(_06927_),
    .Y(_06928_));
 sky130_fd_sc_hd__nand2_1 _14217_ (.A(_06632_),
    .B(_06650_),
    .Y(_06929_));
 sky130_fd_sc_hd__xnor2_1 _14218_ (.A(_06928_),
    .B(_06929_),
    .Y(_06930_));
 sky130_fd_sc_hd__o21ba_1 _14219_ (.A1(_06891_),
    .A2(_06894_),
    .B1_N(_06892_),
    .X(_06931_));
 sky130_fd_sc_hd__xnor2_1 _14220_ (.A(_06930_),
    .B(_06931_),
    .Y(_06932_));
 sky130_fd_sc_hd__o21ai_1 _14221_ (.A1(_06648_),
    .A2(_06645_),
    .B1(_06635_),
    .Y(_06933_));
 sky130_fd_sc_hd__nor3_1 _14222_ (.A(_06860_),
    .B(_06898_),
    .C(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__o21a_1 _14223_ (.A1(_06898_),
    .A2(_06933_),
    .B1(_06860_),
    .X(_06935_));
 sky130_fd_sc_hd__nor2_2 _14224_ (.A(net180),
    .B(_06935_),
    .Y(_06936_));
 sky130_fd_sc_hd__xnor2_1 _14225_ (.A(_06932_),
    .B(_06936_),
    .Y(_06937_));
 sky130_fd_sc_hd__or2b_1 _14226_ (.A(_06895_),
    .B_N(_06896_),
    .X(_06938_));
 sky130_fd_sc_hd__and2b_1 _14227_ (.A_N(_06896_),
    .B(_06895_),
    .X(_06939_));
 sky130_fd_sc_hd__a21oi_1 _14228_ (.A1(_06938_),
    .A2(_06901_),
    .B1(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__nor2_1 _14229_ (.A(_06937_),
    .B(_06940_),
    .Y(_06941_));
 sky130_fd_sc_hd__and2_1 _14230_ (.A(_06937_),
    .B(_06940_),
    .X(_06942_));
 sky130_fd_sc_hd__nor2_1 _14231_ (.A(_06941_),
    .B(_06942_),
    .Y(_06943_));
 sky130_fd_sc_hd__o2bb2a_1 _14232_ (.A1_N(_06632_),
    .A2_N(_06898_),
    .B1(_06899_),
    .B2(_06860_),
    .X(_06944_));
 sky130_fd_sc_hd__nor2_1 _14233_ (.A(_06825_),
    .B(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__and2_1 _14234_ (.A(_06825_),
    .B(_06944_),
    .X(_06946_));
 sky130_fd_sc_hd__nor2_1 _14235_ (.A(_06945_),
    .B(_06946_),
    .Y(_06947_));
 sky130_fd_sc_hd__xnor2_1 _14236_ (.A(_06943_),
    .B(_06947_),
    .Y(_06948_));
 sky130_fd_sc_hd__a21oi_1 _14237_ (.A1(_06905_),
    .A2(_06909_),
    .B1(_06903_),
    .Y(_06949_));
 sky130_fd_sc_hd__nor2_1 _14238_ (.A(_06948_),
    .B(_06949_),
    .Y(_06950_));
 sky130_fd_sc_hd__and2_1 _14239_ (.A(_06948_),
    .B(_06949_),
    .X(_06951_));
 sky130_fd_sc_hd__nor2_1 _14240_ (.A(_06950_),
    .B(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__xnor2_1 _14241_ (.A(_06907_),
    .B(_06952_),
    .Y(_06953_));
 sky130_fd_sc_hd__nor2_1 _14242_ (.A(_06910_),
    .B(_06912_),
    .Y(_06954_));
 sky130_fd_sc_hd__a21oi_1 _14243_ (.A1(_06869_),
    .A2(_06913_),
    .B1(_06954_),
    .Y(_06955_));
 sky130_fd_sc_hd__xnor2_1 _14244_ (.A(_06953_),
    .B(_06955_),
    .Y(_06956_));
 sky130_fd_sc_hd__o21bai_2 _14245_ (.A1(_06919_),
    .A2(_06920_),
    .B1_N(_06917_),
    .Y(_06957_));
 sky130_fd_sc_hd__xnor2_1 _14246_ (.A(_06956_),
    .B(_06957_),
    .Y(_06958_));
 sky130_fd_sc_hd__or2_1 _14247_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[11] ),
    .B(_06168_),
    .X(_06959_));
 sky130_fd_sc_hd__o211a_1 _14248_ (.A1(_06848_),
    .A2(_06958_),
    .B1(_06959_),
    .C1(_06684_),
    .X(_00410_));
 sky130_fd_sc_hd__inv_2 _14249_ (.A(net1090),
    .Y(_06960_));
 sky130_fd_sc_hd__or2b_1 _14250_ (.A(_06931_),
    .B_N(_06930_),
    .X(_06961_));
 sky130_fd_sc_hd__nand2_1 _14251_ (.A(_06932_),
    .B(_06936_),
    .Y(_06962_));
 sky130_fd_sc_hd__inv_2 _14252_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[7] ),
    .Y(_06963_));
 sky130_fd_sc_hd__o2bb2a_1 _14253_ (.A1_N(_06652_),
    .A2_N(\top_inst.grid_inst.data_path_wires[3][6] ),
    .B1(_06630_),
    .B2(_06963_),
    .X(_06964_));
 sky130_fd_sc_hd__and4b_1 _14254_ (.A_N(_06630_),
    .B(\top_inst.grid_inst.data_path_wires[3][6] ),
    .C(_06652_),
    .D(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[7] ),
    .X(_06965_));
 sky130_fd_sc_hd__nand2_1 _14255_ (.A(_06635_),
    .B(_06650_),
    .Y(_06966_));
 sky130_fd_sc_hd__o21a_1 _14256_ (.A1(_06964_),
    .A2(_06965_),
    .B1(_06966_),
    .X(_06967_));
 sky130_fd_sc_hd__nor2_1 _14257_ (.A(_06964_),
    .B(_06965_),
    .Y(_06968_));
 sky130_fd_sc_hd__and3_1 _14258_ (.A(_06635_),
    .B(_06650_),
    .C(_06968_),
    .X(_06969_));
 sky130_fd_sc_hd__nor2_1 _14259_ (.A(_06967_),
    .B(_06969_),
    .Y(_06970_));
 sky130_fd_sc_hd__o21ba_1 _14260_ (.A1(_06926_),
    .A2(_06929_),
    .B1_N(_06927_),
    .X(_06971_));
 sky130_fd_sc_hd__xnor2_1 _14261_ (.A(_06970_),
    .B(_06971_),
    .Y(_06972_));
 sky130_fd_sc_hd__xnor2_1 _14262_ (.A(_06936_),
    .B(_06972_),
    .Y(_06973_));
 sky130_fd_sc_hd__a21o_1 _14263_ (.A1(_06961_),
    .A2(_06962_),
    .B1(_06973_),
    .X(_06974_));
 sky130_fd_sc_hd__nand3_1 _14264_ (.A(_06961_),
    .B(_06962_),
    .C(_06973_),
    .Y(_06975_));
 sky130_fd_sc_hd__nand2_1 _14265_ (.A(_06974_),
    .B(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__o21a_1 _14266_ (.A1(_06640_),
    .A2(_06637_),
    .B1(_06635_),
    .X(_06977_));
 sky130_fd_sc_hd__o21ai_2 _14267_ (.A1(_06898_),
    .A2(net180),
    .B1(_06977_),
    .Y(_06978_));
 sky130_fd_sc_hd__or3_2 _14268_ (.A(_06977_),
    .B(_06898_),
    .C(_06934_),
    .X(_06979_));
 sky130_fd_sc_hd__nand2_2 _14269_ (.A(_06978_),
    .B(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__inv_2 _14270_ (.A(_06980_),
    .Y(_06981_));
 sky130_fd_sc_hd__xnor2_1 _14271_ (.A(_06976_),
    .B(_06981_),
    .Y(_06982_));
 sky130_fd_sc_hd__a21oi_1 _14272_ (.A1(_06943_),
    .A2(_06947_),
    .B1(_06941_),
    .Y(_06983_));
 sky130_fd_sc_hd__xnor2_1 _14273_ (.A(_06982_),
    .B(_06983_),
    .Y(_06984_));
 sky130_fd_sc_hd__xnor2_1 _14274_ (.A(_06945_),
    .B(_06984_),
    .Y(_06985_));
 sky130_fd_sc_hd__a21oi_1 _14275_ (.A1(_06907_),
    .A2(_06952_),
    .B1(_06950_),
    .Y(_06986_));
 sky130_fd_sc_hd__or2_1 _14276_ (.A(_06985_),
    .B(_06986_),
    .X(_06987_));
 sky130_fd_sc_hd__nand2_1 _14277_ (.A(_06985_),
    .B(_06986_),
    .Y(_06988_));
 sky130_fd_sc_hd__nand2_1 _14278_ (.A(_06987_),
    .B(_06988_),
    .Y(_06989_));
 sky130_fd_sc_hd__inv_2 _14279_ (.A(_06956_),
    .Y(_06990_));
 sky130_fd_sc_hd__or2_1 _14280_ (.A(_06953_),
    .B(_06955_),
    .X(_06991_));
 sky130_fd_sc_hd__a21boi_2 _14281_ (.A1(_06990_),
    .A2(_06957_),
    .B1_N(_06991_),
    .Y(_06992_));
 sky130_fd_sc_hd__xnor2_2 _14282_ (.A(_06989_),
    .B(_06992_),
    .Y(_06993_));
 sky130_fd_sc_hd__mux2_1 _14283_ (.A0(_06960_),
    .A1(_06993_),
    .S(_05316_),
    .X(_06994_));
 sky130_fd_sc_hd__nor2_1 _14284_ (.A(_05632_),
    .B(_06994_),
    .Y(_00411_));
 sky130_fd_sc_hd__inv_2 _14285_ (.A(_06978_),
    .Y(_06995_));
 sky130_fd_sc_hd__o21a_1 _14286_ (.A1(_06976_),
    .A2(_06980_),
    .B1(_06974_),
    .X(_06996_));
 sky130_fd_sc_hd__nand2_1 _14287_ (.A(\top_inst.grid_inst.data_path_wires[3][7] ),
    .B(_06652_),
    .Y(_06997_));
 sky130_fd_sc_hd__o21a_1 _14288_ (.A1(_06963_),
    .A2(\top_inst.grid_inst.data_path_wires[3][6] ),
    .B1(_06997_),
    .X(_06998_));
 sky130_fd_sc_hd__nor3_1 _14289_ (.A(_06963_),
    .B(_06632_),
    .C(_06997_),
    .Y(_06999_));
 sky130_fd_sc_hd__nor2_1 _14290_ (.A(_06998_),
    .B(_06999_),
    .Y(_07000_));
 sky130_fd_sc_hd__xnor2_1 _14291_ (.A(_06966_),
    .B(_07000_),
    .Y(_07001_));
 sky130_fd_sc_hd__o21ai_1 _14292_ (.A1(_06965_),
    .A2(_06969_),
    .B1(_07001_),
    .Y(_07002_));
 sky130_fd_sc_hd__or3_1 _14293_ (.A(_06965_),
    .B(_06969_),
    .C(_07001_),
    .X(_07003_));
 sky130_fd_sc_hd__and2_1 _14294_ (.A(_07002_),
    .B(_07003_),
    .X(_07004_));
 sky130_fd_sc_hd__nand2_1 _14295_ (.A(_06936_),
    .B(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__or2_1 _14296_ (.A(_06936_),
    .B(_07004_),
    .X(_07006_));
 sky130_fd_sc_hd__nand2_1 _14297_ (.A(_07005_),
    .B(_07006_),
    .Y(_07007_));
 sky130_fd_sc_hd__or2b_1 _14298_ (.A(_06971_),
    .B_N(_06970_),
    .X(_07008_));
 sky130_fd_sc_hd__a21bo_1 _14299_ (.A1(_06936_),
    .A2(_06972_),
    .B1_N(_07008_),
    .X(_07009_));
 sky130_fd_sc_hd__xor2_1 _14300_ (.A(_07007_),
    .B(_07009_),
    .X(_07010_));
 sky130_fd_sc_hd__xnor2_1 _14301_ (.A(_06981_),
    .B(_07010_),
    .Y(_07011_));
 sky130_fd_sc_hd__and2b_1 _14302_ (.A_N(_06996_),
    .B(_07011_),
    .X(_07012_));
 sky130_fd_sc_hd__and2b_1 _14303_ (.A_N(_07011_),
    .B(_06996_),
    .X(_07013_));
 sky130_fd_sc_hd__nor2_1 _14304_ (.A(_07012_),
    .B(_07013_),
    .Y(_07014_));
 sky130_fd_sc_hd__xnor2_1 _14305_ (.A(_06995_),
    .B(_07014_),
    .Y(_07015_));
 sky130_fd_sc_hd__and2b_1 _14306_ (.A_N(_06983_),
    .B(_06982_),
    .X(_07016_));
 sky130_fd_sc_hd__a21oi_1 _14307_ (.A1(_06945_),
    .A2(_06984_),
    .B1(_07016_),
    .Y(_07017_));
 sky130_fd_sc_hd__nor2_1 _14308_ (.A(_07015_),
    .B(_07017_),
    .Y(_07018_));
 sky130_fd_sc_hd__and2_1 _14309_ (.A(_07015_),
    .B(_07017_),
    .X(_07019_));
 sky130_fd_sc_hd__or2_1 _14310_ (.A(_07018_),
    .B(_07019_),
    .X(_07020_));
 sky130_fd_sc_hd__o21a_1 _14311_ (.A1(_06989_),
    .A2(_06992_),
    .B1(_06987_),
    .X(_07021_));
 sky130_fd_sc_hd__xor2_1 _14312_ (.A(_07020_),
    .B(_07021_),
    .X(_07022_));
 sky130_fd_sc_hd__mux2_1 _14313_ (.A0(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[13] ),
    .A1(_07022_),
    .S(_06701_),
    .X(_07023_));
 sky130_fd_sc_hd__and2_1 _14314_ (.A(_06364_),
    .B(_07023_),
    .X(_07024_));
 sky130_fd_sc_hd__clkbuf_1 _14315_ (.A(_07024_),
    .X(_00412_));
 sky130_fd_sc_hd__or2b_1 _14316_ (.A(_07007_),
    .B_N(_07009_),
    .X(_07025_));
 sky130_fd_sc_hd__o21a_1 _14317_ (.A1(_06980_),
    .A2(_07010_),
    .B1(_07025_),
    .X(_07026_));
 sky130_fd_sc_hd__and3_1 _14318_ (.A(_06635_),
    .B(_06652_),
    .C(_06650_),
    .X(_07027_));
 sky130_fd_sc_hd__o21ba_1 _14319_ (.A1(_06966_),
    .A2(_06998_),
    .B1_N(_06999_),
    .X(_07028_));
 sky130_fd_sc_hd__o211a_1 _14320_ (.A1(_06963_),
    .A2(_06635_),
    .B1(_06966_),
    .C1(_06997_),
    .X(_07029_));
 sky130_fd_sc_hd__o21ba_1 _14321_ (.A1(_07027_),
    .A2(_07028_),
    .B1_N(_07029_),
    .X(_07030_));
 sky130_fd_sc_hd__xnor2_1 _14322_ (.A(_06936_),
    .B(_07030_),
    .Y(_07031_));
 sky130_fd_sc_hd__a21oi_1 _14323_ (.A1(_07002_),
    .A2(_07005_),
    .B1(_07031_),
    .Y(_07032_));
 sky130_fd_sc_hd__and3_1 _14324_ (.A(_07002_),
    .B(_07005_),
    .C(_07031_),
    .X(_07033_));
 sky130_fd_sc_hd__nor2_1 _14325_ (.A(_07032_),
    .B(_07033_),
    .Y(_07034_));
 sky130_fd_sc_hd__xnor2_1 _14326_ (.A(_06980_),
    .B(_07034_),
    .Y(_07035_));
 sky130_fd_sc_hd__and2b_1 _14327_ (.A_N(_07026_),
    .B(_07035_),
    .X(_07036_));
 sky130_fd_sc_hd__and2b_1 _14328_ (.A_N(_07035_),
    .B(_07026_),
    .X(_07037_));
 sky130_fd_sc_hd__nor2_1 _14329_ (.A(_07036_),
    .B(_07037_),
    .Y(_07038_));
 sky130_fd_sc_hd__xnor2_1 _14330_ (.A(_06995_),
    .B(_07038_),
    .Y(_07039_));
 sky130_fd_sc_hd__a21oi_1 _14331_ (.A1(_06995_),
    .A2(_07014_),
    .B1(_07012_),
    .Y(_07040_));
 sky130_fd_sc_hd__or2_1 _14332_ (.A(_07039_),
    .B(_07040_),
    .X(_07041_));
 sky130_fd_sc_hd__nand2_1 _14333_ (.A(_07039_),
    .B(_07040_),
    .Y(_07042_));
 sky130_fd_sc_hd__nand2_1 _14334_ (.A(_07041_),
    .B(_07042_),
    .Y(_07043_));
 sky130_fd_sc_hd__o21ba_1 _14335_ (.A1(_07020_),
    .A2(_07021_),
    .B1_N(_07018_),
    .X(_07044_));
 sky130_fd_sc_hd__nor2_1 _14336_ (.A(_07043_),
    .B(_07044_),
    .Y(_07045_));
 sky130_fd_sc_hd__a21o_1 _14337_ (.A1(_07043_),
    .A2(_07044_),
    .B1(_05633_),
    .X(_07046_));
 sky130_fd_sc_hd__o2bb2a_1 _14338_ (.A1_N(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[14] ),
    .A2_N(_05634_),
    .B1(_07045_),
    .B2(_07046_),
    .X(_07047_));
 sky130_fd_sc_hd__nor2_1 _14339_ (.A(_05632_),
    .B(_07047_),
    .Y(_00413_));
 sky130_fd_sc_hd__buf_4 _14340_ (.A(_05787_),
    .X(_07048_));
 sky130_fd_sc_hd__o21a_1 _14341_ (.A1(_07043_),
    .A2(_07044_),
    .B1(_07041_),
    .X(_07049_));
 sky130_fd_sc_hd__xnor2_2 _14342_ (.A(_06979_),
    .B(_07049_),
    .Y(_07050_));
 sky130_fd_sc_hd__nor2_1 _14343_ (.A(_06936_),
    .B(_07030_),
    .Y(_07051_));
 sky130_fd_sc_hd__a21oi_1 _14344_ (.A1(_06995_),
    .A2(_07038_),
    .B1(_07036_),
    .Y(_07052_));
 sky130_fd_sc_hd__a21oi_1 _14345_ (.A1(_06981_),
    .A2(_07034_),
    .B1(_07032_),
    .Y(_07053_));
 sky130_fd_sc_hd__xnor2_1 _14346_ (.A(_07052_),
    .B(_07053_),
    .Y(_07054_));
 sky130_fd_sc_hd__xnor2_2 _14347_ (.A(_07051_),
    .B(_07054_),
    .Y(_07055_));
 sky130_fd_sc_hd__nor2_1 _14348_ (.A(_07050_),
    .B(_07055_),
    .Y(_07056_));
 sky130_fd_sc_hd__buf_8 _14349_ (.A(_05731_),
    .X(_07057_));
 sky130_fd_sc_hd__a21o_1 _14350_ (.A1(_07050_),
    .A2(_07055_),
    .B1(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__o221a_1 _14351_ (.A1(net1042),
    .A2(_07048_),
    .B1(_07056_),
    .B2(_07058_),
    .C1(_06180_),
    .X(_00414_));
 sky130_fd_sc_hd__buf_8 _14352_ (.A(net34),
    .X(_07059_));
 sky130_fd_sc_hd__mux2_4 _14353_ (.A0(\top_inst.skew_buff_inst.row[1].output_reg[0] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[8] ),
    .S(net206),
    .X(_07060_));
 sky130_fd_sc_hd__clkbuf_4 _14354_ (.A(_07060_),
    .X(_07061_));
 sky130_fd_sc_hd__clkbuf_4 _14355_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[0] ),
    .X(_07062_));
 sky130_fd_sc_hd__or2_1 _14356_ (.A(_07062_),
    .B(_06641_),
    .X(_07063_));
 sky130_fd_sc_hd__o211a_1 _14357_ (.A1(_05290_),
    .A2(_07061_),
    .B1(_07063_),
    .C1(_06684_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_4 _14358_ (.A0(\top_inst.skew_buff_inst.row[1].output_reg[1] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[9] ),
    .S(net208),
    .X(_07064_));
 sky130_fd_sc_hd__buf_4 _14359_ (.A(_07064_),
    .X(_07065_));
 sky130_fd_sc_hd__clkbuf_4 _14360_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[1] ),
    .X(_07066_));
 sky130_fd_sc_hd__or2_1 _14361_ (.A(_07066_),
    .B(_06641_),
    .X(_07067_));
 sky130_fd_sc_hd__o211a_1 _14362_ (.A1(_05290_),
    .A2(_07065_),
    .B1(_07067_),
    .C1(_06684_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_4 _14363_ (.A0(\top_inst.skew_buff_inst.row[1].output_reg[2] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[10] ),
    .S(net187),
    .X(_07068_));
 sky130_fd_sc_hd__buf_6 _14364_ (.A(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__clkbuf_4 _14365_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[2] ),
    .X(_07070_));
 sky130_fd_sc_hd__or2_1 _14366_ (.A(_07070_),
    .B(_06641_),
    .X(_07071_));
 sky130_fd_sc_hd__o211a_1 _14367_ (.A1(_05290_),
    .A2(_07069_),
    .B1(_07071_),
    .C1(_06684_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_4 _14368_ (.A0(\top_inst.skew_buff_inst.row[1].output_reg[3] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[11] ),
    .S(_05266_),
    .X(_07072_));
 sky130_fd_sc_hd__clkbuf_4 _14369_ (.A(_07072_),
    .X(_07073_));
 sky130_fd_sc_hd__buf_2 _14370_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[3] ),
    .X(_07074_));
 sky130_fd_sc_hd__buf_2 _14371_ (.A(_05772_),
    .X(_07075_));
 sky130_fd_sc_hd__or2_1 _14372_ (.A(_07074_),
    .B(_07075_),
    .X(_07076_));
 sky130_fd_sc_hd__o211a_1 _14373_ (.A1(_05290_),
    .A2(_07073_),
    .B1(_07076_),
    .C1(_06684_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_4 _14374_ (.A0(\top_inst.skew_buff_inst.row[1].output_reg[4] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[12] ),
    .S(net207),
    .X(_07077_));
 sky130_fd_sc_hd__clkbuf_4 _14375_ (.A(_07077_),
    .X(_07078_));
 sky130_fd_sc_hd__buf_2 _14376_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[4] ),
    .X(_07079_));
 sky130_fd_sc_hd__or2_1 _14377_ (.A(_07079_),
    .B(_07075_),
    .X(_07080_));
 sky130_fd_sc_hd__o211a_1 _14378_ (.A1(_05290_),
    .A2(_07078_),
    .B1(_07080_),
    .C1(_06684_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_4 _14379_ (.A0(\top_inst.skew_buff_inst.row[1].output_reg[5] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[13] ),
    .S(net208),
    .X(_07081_));
 sky130_fd_sc_hd__buf_2 _14380_ (.A(net1122),
    .X(_07082_));
 sky130_fd_sc_hd__clkbuf_4 _14381_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[5] ),
    .X(_07083_));
 sky130_fd_sc_hd__or2_1 _14382_ (.A(_07083_),
    .B(_07075_),
    .X(_07084_));
 sky130_fd_sc_hd__o211a_1 _14383_ (.A1(_05290_),
    .A2(_07082_),
    .B1(_07084_),
    .C1(_06684_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_4 _14384_ (.A0(\top_inst.skew_buff_inst.row[1].output_reg[6] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[14] ),
    .S(net208),
    .X(_07085_));
 sky130_fd_sc_hd__buf_2 _14385_ (.A(_07085_),
    .X(_07086_));
 sky130_fd_sc_hd__clkbuf_4 _14386_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[6] ),
    .X(_07087_));
 sky130_fd_sc_hd__or2_1 _14387_ (.A(_07087_),
    .B(_07075_),
    .X(_07088_));
 sky130_fd_sc_hd__o211a_1 _14388_ (.A1(_05290_),
    .A2(_07086_),
    .B1(_07088_),
    .C1(_06684_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_2 _14389_ (.A0(\top_inst.skew_buff_inst.row[1].output_reg[7] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[15] ),
    .S(net212),
    .X(_07089_));
 sky130_fd_sc_hd__buf_4 _14390_ (.A(_07089_),
    .X(_07090_));
 sky130_fd_sc_hd__or2_1 _14391_ (.A(_05269_),
    .B(_07090_),
    .X(_07091_));
 sky130_fd_sc_hd__buf_4 _14392_ (.A(_05260_),
    .X(_07092_));
 sky130_fd_sc_hd__o211a_1 _14393_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[7] ),
    .A2(_05276_),
    .B1(_07091_),
    .C1(_07092_),
    .X(_00422_));
 sky130_fd_sc_hd__a21oi_1 _14394_ (.A1(_07062_),
    .A2(_07061_),
    .B1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[0] ),
    .Y(_07093_));
 sky130_fd_sc_hd__and3_1 _14395_ (.A(_07062_),
    .B(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[0] ),
    .C(_07061_),
    .X(_07094_));
 sky130_fd_sc_hd__o21ai_1 _14396_ (.A1(_07093_),
    .A2(_07094_),
    .B1(_05336_),
    .Y(_07095_));
 sky130_fd_sc_hd__o211a_1 _14397_ (.A1(net1077),
    .A2(_06660_),
    .B1(_07095_),
    .C1(_07092_),
    .X(_00423_));
 sky130_fd_sc_hd__a22o_1 _14398_ (.A1(_07066_),
    .A2(_07061_),
    .B1(_07065_),
    .B2(_07062_),
    .X(_07096_));
 sky130_fd_sc_hd__nand4_1 _14399_ (.A(_07066_),
    .B(_07062_),
    .C(_07061_),
    .D(_07065_),
    .Y(_07097_));
 sky130_fd_sc_hd__and3_1 _14400_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[1] ),
    .B(_07096_),
    .C(_07097_),
    .X(_07098_));
 sky130_fd_sc_hd__a21oi_1 _14401_ (.A1(_07096_),
    .A2(_07097_),
    .B1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[1] ),
    .Y(_07099_));
 sky130_fd_sc_hd__o21ba_1 _14402_ (.A1(_07098_),
    .A2(_07099_),
    .B1_N(_07094_),
    .X(_07100_));
 sky130_fd_sc_hd__nor3b_1 _14403_ (.A(_07098_),
    .B(_07099_),
    .C_N(_07094_),
    .Y(_07101_));
 sky130_fd_sc_hd__o21ai_1 _14404_ (.A1(_07100_),
    .A2(_07101_),
    .B1(_05336_),
    .Y(_07102_));
 sky130_fd_sc_hd__o211a_1 _14405_ (.A1(net1045),
    .A2(_06660_),
    .B1(_07102_),
    .C1(_07092_),
    .X(_00424_));
 sky130_fd_sc_hd__a22o_1 _14406_ (.A1(_07066_),
    .A2(_07065_),
    .B1(_07069_),
    .B2(_07062_),
    .X(_07103_));
 sky130_fd_sc_hd__nand4_2 _14407_ (.A(_07066_),
    .B(_07062_),
    .C(_07065_),
    .D(_07069_),
    .Y(_07104_));
 sky130_fd_sc_hd__nand3_1 _14408_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[2] ),
    .B(_07103_),
    .C(_07104_),
    .Y(_07105_));
 sky130_fd_sc_hd__a21o_1 _14409_ (.A1(_07103_),
    .A2(_07104_),
    .B1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[2] ),
    .X(_07106_));
 sky130_fd_sc_hd__nand2_1 _14410_ (.A(_07105_),
    .B(_07106_),
    .Y(_07107_));
 sky130_fd_sc_hd__a21bo_1 _14411_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[1] ),
    .A2(_07096_),
    .B1_N(_07097_),
    .X(_07108_));
 sky130_fd_sc_hd__xnor2_1 _14412_ (.A(_07107_),
    .B(_07108_),
    .Y(_07109_));
 sky130_fd_sc_hd__a21oi_1 _14413_ (.A1(_07070_),
    .A2(_07061_),
    .B1(_07109_),
    .Y(_07110_));
 sky130_fd_sc_hd__and3_1 _14414_ (.A(_07070_),
    .B(_07061_),
    .C(_07109_),
    .X(_07111_));
 sky130_fd_sc_hd__nor2_1 _14415_ (.A(_07110_),
    .B(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__nand2_1 _14416_ (.A(net173),
    .B(_07112_),
    .Y(_07113_));
 sky130_fd_sc_hd__o21a_1 _14417_ (.A1(net173),
    .A2(_07112_),
    .B1(_05315_),
    .X(_07114_));
 sky130_fd_sc_hd__a22o_1 _14418_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[2] ),
    .A2(_06242_),
    .B1(_07113_),
    .B2(_07114_),
    .X(_07115_));
 sky130_fd_sc_hd__and2_1 _14419_ (.A(_06364_),
    .B(_07115_),
    .X(_07116_));
 sky130_fd_sc_hd__clkbuf_1 _14420_ (.A(_07116_),
    .X(_00425_));
 sky130_fd_sc_hd__clkbuf_4 _14421_ (.A(_04869_),
    .X(_07117_));
 sky130_fd_sc_hd__and3_1 _14422_ (.A(_07105_),
    .B(_07106_),
    .C(_07108_),
    .X(_07118_));
 sky130_fd_sc_hd__a22o_1 _14423_ (.A1(_07066_),
    .A2(_07069_),
    .B1(_07073_),
    .B2(_07062_),
    .X(_07119_));
 sky130_fd_sc_hd__nand4_1 _14424_ (.A(_07066_),
    .B(_07062_),
    .C(_07069_),
    .D(_07073_),
    .Y(_07120_));
 sky130_fd_sc_hd__and3_1 _14425_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[3] ),
    .B(_07119_),
    .C(_07120_),
    .X(_07121_));
 sky130_fd_sc_hd__a21oi_1 _14426_ (.A1(_07119_),
    .A2(_07120_),
    .B1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[3] ),
    .Y(_07122_));
 sky130_fd_sc_hd__a211oi_1 _14427_ (.A1(_07104_),
    .A2(_07105_),
    .B1(_07121_),
    .C1(_07122_),
    .Y(_07123_));
 sky130_fd_sc_hd__o211ai_1 _14428_ (.A1(_07121_),
    .A2(_07122_),
    .B1(_07104_),
    .C1(_07105_),
    .Y(_07124_));
 sky130_fd_sc_hd__or2b_1 _14429_ (.A(_07123_),
    .B_N(_07124_),
    .X(_07125_));
 sky130_fd_sc_hd__a22o_1 _14430_ (.A1(_07074_),
    .A2(_07061_),
    .B1(_07065_),
    .B2(_07070_),
    .X(_07126_));
 sky130_fd_sc_hd__nand4_2 _14431_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[3] ),
    .B(_07070_),
    .C(_07060_),
    .D(_07065_),
    .Y(_07127_));
 sky130_fd_sc_hd__nand2_1 _14432_ (.A(_07126_),
    .B(_07127_),
    .Y(_07128_));
 sky130_fd_sc_hd__xor2_1 _14433_ (.A(_07125_),
    .B(_07128_),
    .X(_07129_));
 sky130_fd_sc_hd__o21a_1 _14434_ (.A1(_07118_),
    .A2(_07111_),
    .B1(_07129_),
    .X(_07130_));
 sky130_fd_sc_hd__or3_1 _14435_ (.A(_07118_),
    .B(_07111_),
    .C(_07129_),
    .X(_07131_));
 sky130_fd_sc_hd__and2b_1 _14436_ (.A_N(_07130_),
    .B(_07131_),
    .X(_07132_));
 sky130_fd_sc_hd__xnor2_1 _14437_ (.A(_07113_),
    .B(_07132_),
    .Y(_07133_));
 sky130_fd_sc_hd__mux2_1 _14438_ (.A0(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[3] ),
    .A1(_07133_),
    .S(_06701_),
    .X(_07134_));
 sky130_fd_sc_hd__and2_1 _14439_ (.A(_07117_),
    .B(_07134_),
    .X(_07135_));
 sky130_fd_sc_hd__clkbuf_1 _14440_ (.A(_07135_),
    .X(_00426_));
 sky130_fd_sc_hd__a22o_1 _14441_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[1] ),
    .A2(_07072_),
    .B1(_07077_),
    .B2(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[0] ),
    .X(_07136_));
 sky130_fd_sc_hd__nand4_1 _14442_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[1] ),
    .B(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[0] ),
    .C(_07072_),
    .D(_07077_),
    .Y(_07137_));
 sky130_fd_sc_hd__and3_1 _14443_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[4] ),
    .B(_07136_),
    .C(_07137_),
    .X(_07138_));
 sky130_fd_sc_hd__a21oi_1 _14444_ (.A1(_07136_),
    .A2(_07137_),
    .B1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[4] ),
    .Y(_07139_));
 sky130_fd_sc_hd__or3_1 _14445_ (.A(_07127_),
    .B(_07138_),
    .C(_07139_),
    .X(_07140_));
 sky130_fd_sc_hd__o21ai_1 _14446_ (.A1(_07138_),
    .A2(_07139_),
    .B1(_07127_),
    .Y(_07141_));
 sky130_fd_sc_hd__a21bo_1 _14447_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[3] ),
    .A2(_07119_),
    .B1_N(_07120_),
    .X(_07142_));
 sky130_fd_sc_hd__nand3_1 _14448_ (.A(_07140_),
    .B(_07141_),
    .C(_07142_),
    .Y(_07143_));
 sky130_fd_sc_hd__a21o_1 _14449_ (.A1(_07140_),
    .A2(_07141_),
    .B1(_07142_),
    .X(_07144_));
 sky130_fd_sc_hd__nand2_1 _14450_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[2] ),
    .B(_07069_),
    .Y(_07145_));
 sky130_fd_sc_hd__nand4_4 _14451_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[3] ),
    .C(_07060_),
    .D(_07064_),
    .Y(_07146_));
 sky130_fd_sc_hd__a22o_1 _14452_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[4] ),
    .A2(_07060_),
    .B1(_07064_),
    .B2(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[3] ),
    .X(_07147_));
 sky130_fd_sc_hd__nand3b_2 _14453_ (.A_N(_07145_),
    .B(_07146_),
    .C(_07147_),
    .Y(_07148_));
 sky130_fd_sc_hd__a21bo_1 _14454_ (.A1(_07146_),
    .A2(_07147_),
    .B1_N(_07145_),
    .X(_07149_));
 sky130_fd_sc_hd__and2_1 _14455_ (.A(_07148_),
    .B(_07149_),
    .X(_07150_));
 sky130_fd_sc_hd__and3_1 _14456_ (.A(_07143_),
    .B(_07144_),
    .C(_07150_),
    .X(_07151_));
 sky130_fd_sc_hd__a21oi_1 _14457_ (.A1(_07143_),
    .A2(_07144_),
    .B1(_07150_),
    .Y(_07152_));
 sky130_fd_sc_hd__a31o_1 _14458_ (.A1(_07124_),
    .A2(_07126_),
    .A3(_07127_),
    .B1(_07123_),
    .X(_07153_));
 sky130_fd_sc_hd__or3b_2 _14459_ (.A(net1125),
    .B(_07152_),
    .C_N(_07153_),
    .X(_07154_));
 sky130_fd_sc_hd__o21bai_2 _14460_ (.A1(net1125),
    .A2(_07152_),
    .B1_N(_07153_),
    .Y(_07155_));
 sky130_fd_sc_hd__nand2_1 _14461_ (.A(_07154_),
    .B(_07155_),
    .Y(_07156_));
 sky130_fd_sc_hd__a31o_1 _14462_ (.A1(net173),
    .A2(_07112_),
    .A3(_07131_),
    .B1(_07130_),
    .X(_07157_));
 sky130_fd_sc_hd__nor2_1 _14463_ (.A(_07156_),
    .B(_07157_),
    .Y(_07158_));
 sky130_fd_sc_hd__a21o_1 _14464_ (.A1(_07156_),
    .A2(_07157_),
    .B1(_07057_),
    .X(_07159_));
 sky130_fd_sc_hd__o221a_1 _14465_ (.A1(net1070),
    .A2(_07048_),
    .B1(_07158_),
    .B2(_07159_),
    .C1(_06180_),
    .X(_00427_));
 sky130_fd_sc_hd__inv_2 _14466_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[5] ),
    .Y(_07160_));
 sky130_fd_sc_hd__and4b_1 _14467_ (.A_N(_07113_),
    .B(_07132_),
    .C(_07154_),
    .D(_07155_),
    .X(_07161_));
 sky130_fd_sc_hd__a21bo_1 _14468_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[4] ),
    .A2(_07136_),
    .B1_N(_07137_),
    .X(_07162_));
 sky130_fd_sc_hd__a22o_1 _14469_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[1] ),
    .A2(_07077_),
    .B1(_07081_),
    .B2(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[0] ),
    .X(_07163_));
 sky130_fd_sc_hd__nand4_1 _14470_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[1] ),
    .B(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[0] ),
    .C(_07077_),
    .D(_07081_),
    .Y(_07164_));
 sky130_fd_sc_hd__and3_1 _14471_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[5] ),
    .B(_07163_),
    .C(_07164_),
    .X(_07165_));
 sky130_fd_sc_hd__a21oi_1 _14472_ (.A1(_07163_),
    .A2(_07164_),
    .B1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[5] ),
    .Y(_07166_));
 sky130_fd_sc_hd__a211o_1 _14473_ (.A1(_07146_),
    .A2(_07148_),
    .B1(_07165_),
    .C1(_07166_),
    .X(_07167_));
 sky130_fd_sc_hd__o211ai_2 _14474_ (.A1(_07165_),
    .A2(_07166_),
    .B1(_07146_),
    .C1(_07148_),
    .Y(_07168_));
 sky130_fd_sc_hd__nand3_2 _14475_ (.A(_07162_),
    .B(_07167_),
    .C(_07168_),
    .Y(_07169_));
 sky130_fd_sc_hd__a21o_1 _14476_ (.A1(_07167_),
    .A2(_07168_),
    .B1(_07162_),
    .X(_07170_));
 sky130_fd_sc_hd__a22o_1 _14477_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[4] ),
    .A2(_07064_),
    .B1(_07068_),
    .B2(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[3] ),
    .X(_07171_));
 sky130_fd_sc_hd__nand4_4 _14478_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[3] ),
    .C(_07064_),
    .D(_07068_),
    .Y(_07172_));
 sky130_fd_sc_hd__nand4_2 _14479_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[2] ),
    .B(_07073_),
    .C(_07171_),
    .D(_07172_),
    .Y(_07173_));
 sky130_fd_sc_hd__a22o_1 _14480_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[2] ),
    .A2(_07073_),
    .B1(_07171_),
    .B2(_07172_),
    .X(_07174_));
 sky130_fd_sc_hd__and4_1 _14481_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[5] ),
    .B(_07060_),
    .C(_07173_),
    .D(_07174_),
    .X(_07175_));
 sky130_fd_sc_hd__a22oi_1 _14482_ (.A1(_07083_),
    .A2(_07061_),
    .B1(_07173_),
    .B2(_07174_),
    .Y(_07176_));
 sky130_fd_sc_hd__nor2_1 _14483_ (.A(_07175_),
    .B(_07176_),
    .Y(_07177_));
 sky130_fd_sc_hd__and3_1 _14484_ (.A(_07169_),
    .B(_07170_),
    .C(_07177_),
    .X(_07178_));
 sky130_fd_sc_hd__a21oi_1 _14485_ (.A1(_07169_),
    .A2(_07170_),
    .B1(_07177_),
    .Y(_07179_));
 sky130_fd_sc_hd__nor3b_2 _14486_ (.A(_07178_),
    .B(_07179_),
    .C_N(_07151_),
    .Y(_07180_));
 sky130_fd_sc_hd__o21ba_1 _14487_ (.A1(_07178_),
    .A2(_07179_),
    .B1_N(net1125),
    .X(_07181_));
 sky130_fd_sc_hd__nand2_1 _14488_ (.A(_07140_),
    .B(_07143_),
    .Y(_07182_));
 sky130_fd_sc_hd__nor3b_1 _14489_ (.A(net171),
    .B(_07181_),
    .C_N(_07182_),
    .Y(_07183_));
 sky130_fd_sc_hd__o21ba_1 _14490_ (.A1(_07180_),
    .A2(_07181_),
    .B1_N(_07182_),
    .X(_07184_));
 sky130_fd_sc_hd__or2_2 _14491_ (.A(_07183_),
    .B(_07184_),
    .X(_07185_));
 sky130_fd_sc_hd__nor3b_1 _14492_ (.A(net1125),
    .B(_07152_),
    .C_N(_07153_),
    .Y(_07186_));
 sky130_fd_sc_hd__a21o_1 _14493_ (.A1(_07130_),
    .A2(_07155_),
    .B1(_07186_),
    .X(_07187_));
 sky130_fd_sc_hd__xnor2_1 _14494_ (.A(_07185_),
    .B(_07187_),
    .Y(_07188_));
 sky130_fd_sc_hd__xnor2_1 _14495_ (.A(_07161_),
    .B(_07188_),
    .Y(_07189_));
 sky130_fd_sc_hd__mux2_1 _14496_ (.A0(_07160_),
    .A1(_07189_),
    .S(_05316_),
    .X(_07190_));
 sky130_fd_sc_hd__nor2_1 _14497_ (.A(_05632_),
    .B(_07190_),
    .Y(_00428_));
 sky130_fd_sc_hd__a21bo_1 _14498_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[5] ),
    .A2(_07163_),
    .B1_N(_07164_),
    .X(_07191_));
 sky130_fd_sc_hd__a22o_1 _14499_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[1] ),
    .A2(_07081_),
    .B1(_07085_),
    .B2(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[0] ),
    .X(_07192_));
 sky130_fd_sc_hd__nand4_1 _14500_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[1] ),
    .B(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[0] ),
    .C(_07081_),
    .D(_07085_),
    .Y(_07193_));
 sky130_fd_sc_hd__and3_1 _14501_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[6] ),
    .B(_07192_),
    .C(_07193_),
    .X(_07194_));
 sky130_fd_sc_hd__a21oi_1 _14502_ (.A1(_07192_),
    .A2(_07193_),
    .B1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[6] ),
    .Y(_07195_));
 sky130_fd_sc_hd__a211o_1 _14503_ (.A1(_07172_),
    .A2(_07173_),
    .B1(_07194_),
    .C1(_07195_),
    .X(_07196_));
 sky130_fd_sc_hd__o211ai_2 _14504_ (.A1(_07194_),
    .A2(_07195_),
    .B1(_07172_),
    .C1(_07173_),
    .Y(_07197_));
 sky130_fd_sc_hd__nand3_2 _14505_ (.A(_07191_),
    .B(_07196_),
    .C(_07197_),
    .Y(_07198_));
 sky130_fd_sc_hd__a21o_1 _14506_ (.A1(_07196_),
    .A2(_07197_),
    .B1(_07191_),
    .X(_07199_));
 sky130_fd_sc_hd__nand4_2 _14507_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[3] ),
    .C(_07068_),
    .D(_07072_),
    .Y(_07200_));
 sky130_fd_sc_hd__a22o_1 _14508_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[4] ),
    .A2(_07068_),
    .B1(_07072_),
    .B2(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[3] ),
    .X(_07201_));
 sky130_fd_sc_hd__nand4_2 _14509_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[2] ),
    .B(_07078_),
    .C(_07200_),
    .D(_07201_),
    .Y(_07202_));
 sky130_fd_sc_hd__a22o_1 _14510_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[2] ),
    .A2(_07078_),
    .B1(_07200_),
    .B2(_07201_),
    .X(_07203_));
 sky130_fd_sc_hd__a22oi_1 _14511_ (.A1(_07087_),
    .A2(_07060_),
    .B1(_07065_),
    .B2(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[5] ),
    .Y(_07204_));
 sky130_fd_sc_hd__and4_1 _14512_ (.A(_07087_),
    .B(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[5] ),
    .C(_07060_),
    .D(_07065_),
    .X(_07205_));
 sky130_fd_sc_hd__nor2_1 _14513_ (.A(_07204_),
    .B(_07205_),
    .Y(_07206_));
 sky130_fd_sc_hd__nand3_1 _14514_ (.A(_07202_),
    .B(_07203_),
    .C(_07206_),
    .Y(_07207_));
 sky130_fd_sc_hd__a21o_1 _14515_ (.A1(_07202_),
    .A2(_07203_),
    .B1(_07206_),
    .X(_07208_));
 sky130_fd_sc_hd__nand3_1 _14516_ (.A(_07175_),
    .B(_07207_),
    .C(_07208_),
    .Y(_07209_));
 sky130_fd_sc_hd__a21o_1 _14517_ (.A1(_07207_),
    .A2(_07208_),
    .B1(_07175_),
    .X(_07210_));
 sky130_fd_sc_hd__nand4_1 _14518_ (.A(_07198_),
    .B(_07199_),
    .C(_07209_),
    .D(_07210_),
    .Y(_07211_));
 sky130_fd_sc_hd__a22o_1 _14519_ (.A1(_07198_),
    .A2(_07199_),
    .B1(_07209_),
    .B2(_07210_),
    .X(_07212_));
 sky130_fd_sc_hd__and3_1 _14520_ (.A(_07178_),
    .B(_07211_),
    .C(_07212_),
    .X(_07213_));
 sky130_fd_sc_hd__a21oi_1 _14521_ (.A1(_07211_),
    .A2(_07212_),
    .B1(_07178_),
    .Y(_07214_));
 sky130_fd_sc_hd__a211o_1 _14522_ (.A1(net209),
    .A2(_07169_),
    .B1(_07213_),
    .C1(_07214_),
    .X(_07215_));
 sky130_fd_sc_hd__o211ai_1 _14523_ (.A1(_07213_),
    .A2(_07214_),
    .B1(net209),
    .C1(_07169_),
    .Y(_07216_));
 sky130_fd_sc_hd__o211a_1 _14524_ (.A1(net171),
    .A2(_07183_),
    .B1(_07215_),
    .C1(_07216_),
    .X(_07217_));
 sky130_fd_sc_hd__a211oi_1 _14525_ (.A1(_07215_),
    .A2(_07216_),
    .B1(net171),
    .C1(_07183_),
    .Y(_07218_));
 sky130_fd_sc_hd__nor4_4 _14526_ (.A(_07154_),
    .B(_07185_),
    .C(_07217_),
    .D(_07218_),
    .Y(_07219_));
 sky130_fd_sc_hd__o22a_1 _14527_ (.A1(_07154_),
    .A2(_07185_),
    .B1(_07217_),
    .B2(_07218_),
    .X(_07220_));
 sky130_fd_sc_hd__nor2_1 _14528_ (.A(_07219_),
    .B(_07220_),
    .Y(_07221_));
 sky130_fd_sc_hd__nand3_1 _14529_ (.A(_07130_),
    .B(_07154_),
    .C(_07155_),
    .Y(_07222_));
 sky130_fd_sc_hd__a2bb2o_2 _14530_ (.A1_N(_07185_),
    .A2_N(_07222_),
    .B1(_07188_),
    .B2(_07161_),
    .X(_07223_));
 sky130_fd_sc_hd__xor2_1 _14531_ (.A(_07221_),
    .B(_07223_),
    .X(_07224_));
 sky130_fd_sc_hd__mux2_1 _14532_ (.A0(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[6] ),
    .A1(_07224_),
    .S(_06701_),
    .X(_07225_));
 sky130_fd_sc_hd__and2_1 _14533_ (.A(_07117_),
    .B(_07225_),
    .X(_07226_));
 sky130_fd_sc_hd__clkbuf_1 _14534_ (.A(_07226_),
    .X(_00429_));
 sky130_fd_sc_hd__a21boi_2 _14535_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[6] ),
    .A2(_07192_),
    .B1_N(_07193_),
    .Y(_07227_));
 sky130_fd_sc_hd__nand2_1 _14536_ (.A(_07200_),
    .B(_07202_),
    .Y(_07228_));
 sky130_fd_sc_hd__and3_1 _14537_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[0] ),
    .B(_07085_),
    .C(_07089_),
    .X(_07229_));
 sky130_fd_sc_hd__a22o_1 _14538_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[1] ),
    .A2(_07085_),
    .B1(_07089_),
    .B2(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[0] ),
    .X(_07230_));
 sky130_fd_sc_hd__a21bo_1 _14539_ (.A1(_07066_),
    .A2(_07229_),
    .B1_N(_07230_),
    .X(_07231_));
 sky130_fd_sc_hd__xor2_1 _14540_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[7] ),
    .B(_07231_),
    .X(_07232_));
 sky130_fd_sc_hd__xnor2_1 _14541_ (.A(_07228_),
    .B(_07232_),
    .Y(_07233_));
 sky130_fd_sc_hd__xnor2_1 _14542_ (.A(_07227_),
    .B(_07233_),
    .Y(_07234_));
 sky130_fd_sc_hd__and3_1 _14543_ (.A(_07202_),
    .B(_07203_),
    .C(_07206_),
    .X(_07235_));
 sky130_fd_sc_hd__nand2_1 _14544_ (.A(_07070_),
    .B(_07081_),
    .Y(_07236_));
 sky130_fd_sc_hd__a22oi_1 _14545_ (.A1(_07079_),
    .A2(_07073_),
    .B1(_07077_),
    .B2(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[3] ),
    .Y(_07237_));
 sky130_fd_sc_hd__and4_1 _14546_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[3] ),
    .C(_07072_),
    .D(_07077_),
    .X(_07238_));
 sky130_fd_sc_hd__nor2_1 _14547_ (.A(_07237_),
    .B(_07238_),
    .Y(_07239_));
 sky130_fd_sc_hd__xnor2_1 _14548_ (.A(_07236_),
    .B(_07239_),
    .Y(_07240_));
 sky130_fd_sc_hd__inv_2 _14549_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[7] ),
    .Y(_07241_));
 sky130_fd_sc_hd__inv_2 _14550_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[6] ),
    .Y(_07242_));
 sky130_fd_sc_hd__or4b_4 _14551_ (.A(_07241_),
    .B(_07242_),
    .C(_07060_),
    .D_N(_07064_),
    .X(_07243_));
 sky130_fd_sc_hd__a2bb2o_1 _14552_ (.A1_N(_07241_),
    .A2_N(_07060_),
    .B1(_07064_),
    .B2(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[6] ),
    .X(_07244_));
 sky130_fd_sc_hd__nand4_1 _14553_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[5] ),
    .B(_07069_),
    .C(_07243_),
    .D(_07244_),
    .Y(_07245_));
 sky130_fd_sc_hd__a22o_1 _14554_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[5] ),
    .A2(_07069_),
    .B1(_07243_),
    .B2(_07244_),
    .X(_07246_));
 sky130_fd_sc_hd__nand3_1 _14555_ (.A(_07205_),
    .B(_07245_),
    .C(_07246_),
    .Y(_07247_));
 sky130_fd_sc_hd__a21o_1 _14556_ (.A1(_07245_),
    .A2(_07246_),
    .B1(_07205_),
    .X(_07248_));
 sky130_fd_sc_hd__nand3_1 _14557_ (.A(_07240_),
    .B(_07247_),
    .C(_07248_),
    .Y(_07249_));
 sky130_fd_sc_hd__a21o_1 _14558_ (.A1(_07247_),
    .A2(_07248_),
    .B1(_07240_),
    .X(_07250_));
 sky130_fd_sc_hd__nand3_1 _14559_ (.A(_07235_),
    .B(_07249_),
    .C(_07250_),
    .Y(_07251_));
 sky130_fd_sc_hd__a21o_1 _14560_ (.A1(_07249_),
    .A2(_07250_),
    .B1(_07235_),
    .X(_07252_));
 sky130_fd_sc_hd__nand3_1 _14561_ (.A(_07234_),
    .B(_07251_),
    .C(_07252_),
    .Y(_07253_));
 sky130_fd_sc_hd__a21o_1 _14562_ (.A1(_07251_),
    .A2(_07252_),
    .B1(_07234_),
    .X(_07254_));
 sky130_fd_sc_hd__nand2_1 _14563_ (.A(_07209_),
    .B(_07211_),
    .Y(_07255_));
 sky130_fd_sc_hd__and3_1 _14564_ (.A(_07253_),
    .B(_07254_),
    .C(_07255_),
    .X(_07256_));
 sky130_fd_sc_hd__a21oi_1 _14565_ (.A1(_07253_),
    .A2(_07254_),
    .B1(_07255_),
    .Y(_07257_));
 sky130_fd_sc_hd__a211oi_1 _14566_ (.A1(net230),
    .A2(_07198_),
    .B1(_07256_),
    .C1(_07257_),
    .Y(_07258_));
 sky130_fd_sc_hd__o211a_1 _14567_ (.A1(_07256_),
    .A2(_07257_),
    .B1(net230),
    .C1(_07198_),
    .X(_07259_));
 sky130_fd_sc_hd__and2b_1 _14568_ (.A_N(_07213_),
    .B(_07215_),
    .X(_07260_));
 sky130_fd_sc_hd__or3_4 _14569_ (.A(_07258_),
    .B(_07259_),
    .C(_07260_),
    .X(_07261_));
 sky130_fd_sc_hd__o21ai_1 _14570_ (.A1(_07258_),
    .A2(_07259_),
    .B1(_07260_),
    .Y(_07262_));
 sky130_fd_sc_hd__nand3_1 _14571_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[7] ),
    .B(_07261_),
    .C(_07262_),
    .Y(_07263_));
 sky130_fd_sc_hd__a21o_1 _14572_ (.A1(_07261_),
    .A2(_07262_),
    .B1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[7] ),
    .X(_07264_));
 sky130_fd_sc_hd__and3_1 _14573_ (.A(_07217_),
    .B(_07263_),
    .C(_07264_),
    .X(_07265_));
 sky130_fd_sc_hd__a21oi_1 _14574_ (.A1(_07263_),
    .A2(_07264_),
    .B1(_07217_),
    .Y(_07266_));
 sky130_fd_sc_hd__nor2_1 _14575_ (.A(_07265_),
    .B(_07266_),
    .Y(_07267_));
 sky130_fd_sc_hd__a21oi_2 _14576_ (.A1(_07221_),
    .A2(_07223_),
    .B1(_07219_),
    .Y(_07268_));
 sky130_fd_sc_hd__xnor2_1 _14577_ (.A(_07267_),
    .B(_07268_),
    .Y(_07269_));
 sky130_fd_sc_hd__mux2_1 _14578_ (.A0(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[7] ),
    .A1(_07269_),
    .S(_06701_),
    .X(_07270_));
 sky130_fd_sc_hd__and2_1 _14579_ (.A(_07117_),
    .B(_07270_),
    .X(_07271_));
 sky130_fd_sc_hd__clkbuf_1 _14580_ (.A(_07271_),
    .X(_00430_));
 sky130_fd_sc_hd__or2_1 _14581_ (.A(_07256_),
    .B(_07258_),
    .X(_07272_));
 sky130_fd_sc_hd__or2b_1 _14582_ (.A(_07232_),
    .B_N(_07228_),
    .X(_07273_));
 sky130_fd_sc_hd__or2b_1 _14583_ (.A(_07227_),
    .B_N(_07233_),
    .X(_07274_));
 sky130_fd_sc_hd__nand2_1 _14584_ (.A(_07273_),
    .B(_07274_),
    .Y(_07275_));
 sky130_fd_sc_hd__a22o_1 _14585_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[7] ),
    .A2(_07230_),
    .B1(_07229_),
    .B2(_07066_),
    .X(_07276_));
 sky130_fd_sc_hd__a31o_1 _14586_ (.A1(_07070_),
    .A2(_07082_),
    .A3(_07239_),
    .B1(_07238_),
    .X(_07277_));
 sky130_fd_sc_hd__o21ai_2 _14587_ (.A1(_07066_),
    .A2(_07062_),
    .B1(_07090_),
    .Y(_07278_));
 sky130_fd_sc_hd__and3_1 _14588_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[1] ),
    .B(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[0] ),
    .C(_07089_),
    .X(_07279_));
 sky130_fd_sc_hd__clkbuf_4 _14589_ (.A(_07279_),
    .X(_07280_));
 sky130_fd_sc_hd__nor2_4 _14590_ (.A(_07278_),
    .B(_07280_),
    .Y(_07281_));
 sky130_fd_sc_hd__xnor2_1 _14591_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[8] ),
    .B(_07281_),
    .Y(_07282_));
 sky130_fd_sc_hd__xnor2_1 _14592_ (.A(_07277_),
    .B(_07282_),
    .Y(_07283_));
 sky130_fd_sc_hd__xor2_1 _14593_ (.A(_07276_),
    .B(_07283_),
    .X(_07284_));
 sky130_fd_sc_hd__nand2_1 _14594_ (.A(_07070_),
    .B(_07086_),
    .Y(_07285_));
 sky130_fd_sc_hd__a22oi_1 _14595_ (.A1(_07079_),
    .A2(_07078_),
    .B1(_07082_),
    .B2(_07074_),
    .Y(_07286_));
 sky130_fd_sc_hd__and4_1 _14596_ (.A(_07079_),
    .B(_07074_),
    .C(_07078_),
    .D(_07082_),
    .X(_07287_));
 sky130_fd_sc_hd__nor2_1 _14597_ (.A(_07286_),
    .B(_07287_),
    .Y(_07288_));
 sky130_fd_sc_hd__xnor2_2 _14598_ (.A(_07285_),
    .B(_07288_),
    .Y(_07289_));
 sky130_fd_sc_hd__inv_2 _14599_ (.A(_07068_),
    .Y(_07290_));
 sky130_fd_sc_hd__or4_4 _14600_ (.A(_07241_),
    .B(_07242_),
    .C(_07065_),
    .D(_07290_),
    .X(_07291_));
 sky130_fd_sc_hd__inv_2 _14601_ (.A(_07064_),
    .Y(_07292_));
 sky130_fd_sc_hd__a22o_1 _14602_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[7] ),
    .A2(_07292_),
    .B1(_07069_),
    .B2(_07087_),
    .X(_07293_));
 sky130_fd_sc_hd__nand4_1 _14603_ (.A(_07083_),
    .B(_07073_),
    .C(_07291_),
    .D(_07293_),
    .Y(_07294_));
 sky130_fd_sc_hd__a22o_1 _14604_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[5] ),
    .A2(_07073_),
    .B1(_07291_),
    .B2(_07293_),
    .X(_07295_));
 sky130_fd_sc_hd__nand2_2 _14605_ (.A(_07294_),
    .B(_07295_),
    .Y(_07296_));
 sky130_fd_sc_hd__and2_1 _14606_ (.A(_07243_),
    .B(_07245_),
    .X(_07297_));
 sky130_fd_sc_hd__xor2_2 _14607_ (.A(_07296_),
    .B(_07297_),
    .X(_07298_));
 sky130_fd_sc_hd__xnor2_2 _14608_ (.A(_07289_),
    .B(_07298_),
    .Y(_07299_));
 sky130_fd_sc_hd__and2_1 _14609_ (.A(_07247_),
    .B(_07249_),
    .X(_07300_));
 sky130_fd_sc_hd__xor2_1 _14610_ (.A(_07299_),
    .B(_07300_),
    .X(_07301_));
 sky130_fd_sc_hd__xnor2_1 _14611_ (.A(_07284_),
    .B(_07301_),
    .Y(_07302_));
 sky130_fd_sc_hd__nand2_1 _14612_ (.A(_07251_),
    .B(_07253_),
    .Y(_07303_));
 sky130_fd_sc_hd__xor2_1 _14613_ (.A(_07302_),
    .B(_07303_),
    .X(_07304_));
 sky130_fd_sc_hd__xnor2_1 _14614_ (.A(_07275_),
    .B(_07304_),
    .Y(_07305_));
 sky130_fd_sc_hd__xnor2_1 _14615_ (.A(_07272_),
    .B(_07305_),
    .Y(_07306_));
 sky130_fd_sc_hd__nand2_1 _14616_ (.A(_07261_),
    .B(_07263_),
    .Y(_07307_));
 sky130_fd_sc_hd__xnor2_1 _14617_ (.A(_07306_),
    .B(_07307_),
    .Y(_07308_));
 sky130_fd_sc_hd__o21bai_2 _14618_ (.A1(_07266_),
    .A2(_07268_),
    .B1_N(_07265_),
    .Y(_07309_));
 sky130_fd_sc_hd__and2_1 _14619_ (.A(_07308_),
    .B(_07309_),
    .X(_07310_));
 sky130_fd_sc_hd__o21ai_1 _14620_ (.A1(_07308_),
    .A2(_07309_),
    .B1(_05335_),
    .Y(_07311_));
 sky130_fd_sc_hd__o2bb2a_1 _14621_ (.A1_N(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[8] ),
    .A2_N(_05634_),
    .B1(_07310_),
    .B2(_07311_),
    .X(_07312_));
 sky130_fd_sc_hd__nor2_1 _14622_ (.A(_05632_),
    .B(_07312_),
    .Y(_00431_));
 sky130_fd_sc_hd__nand2_1 _14623_ (.A(_07272_),
    .B(_07305_),
    .Y(_07313_));
 sky130_fd_sc_hd__inv_2 _14624_ (.A(_07313_),
    .Y(_07314_));
 sky130_fd_sc_hd__and2b_1 _14625_ (.A_N(_07306_),
    .B(_07307_),
    .X(_07315_));
 sky130_fd_sc_hd__a21o_1 _14626_ (.A1(_07308_),
    .A2(_07309_),
    .B1(_07315_),
    .X(_07316_));
 sky130_fd_sc_hd__or2b_1 _14627_ (.A(_07282_),
    .B_N(_07277_),
    .X(_07317_));
 sky130_fd_sc_hd__a21bo_2 _14628_ (.A1(_07276_),
    .A2(_07283_),
    .B1_N(_07317_),
    .X(_07318_));
 sky130_fd_sc_hd__a21oi_1 _14629_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[8] ),
    .A2(_07281_),
    .B1(_07280_),
    .Y(_07319_));
 sky130_fd_sc_hd__xnor2_1 _14630_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[9] ),
    .B(_07281_),
    .Y(_07320_));
 sky130_fd_sc_hd__a31o_1 _14631_ (.A1(_07070_),
    .A2(_07086_),
    .A3(_07288_),
    .B1(_07287_),
    .X(_07321_));
 sky130_fd_sc_hd__and2b_1 _14632_ (.A_N(_07320_),
    .B(_07321_),
    .X(_07322_));
 sky130_fd_sc_hd__and2b_1 _14633_ (.A_N(_07321_),
    .B(_07320_),
    .X(_07323_));
 sky130_fd_sc_hd__nor2_1 _14634_ (.A(_07322_),
    .B(_07323_),
    .Y(_07324_));
 sky130_fd_sc_hd__xnor2_1 _14635_ (.A(_07319_),
    .B(_07324_),
    .Y(_07325_));
 sky130_fd_sc_hd__nor2_1 _14636_ (.A(_07296_),
    .B(_07297_),
    .Y(_07326_));
 sky130_fd_sc_hd__and2_1 _14637_ (.A(_07289_),
    .B(_07298_),
    .X(_07327_));
 sky130_fd_sc_hd__nand2_4 _14638_ (.A(_07070_),
    .B(_07090_),
    .Y(_07328_));
 sky130_fd_sc_hd__a22o_1 _14639_ (.A1(_07079_),
    .A2(_07082_),
    .B1(_07086_),
    .B2(_07074_),
    .X(_07329_));
 sky130_fd_sc_hd__nand4_1 _14640_ (.A(_07079_),
    .B(_07074_),
    .C(_07082_),
    .D(_07086_),
    .Y(_07330_));
 sky130_fd_sc_hd__nand2_1 _14641_ (.A(_07329_),
    .B(_07330_),
    .Y(_07331_));
 sky130_fd_sc_hd__xor2_1 _14642_ (.A(_07328_),
    .B(_07331_),
    .X(_07332_));
 sky130_fd_sc_hd__inv_2 _14643_ (.A(_07072_),
    .Y(_07333_));
 sky130_fd_sc_hd__or4_4 _14644_ (.A(_07241_),
    .B(_07242_),
    .C(_07069_),
    .D(_07333_),
    .X(_07334_));
 sky130_fd_sc_hd__a22o_1 _14645_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[7] ),
    .A2(_07290_),
    .B1(_07073_),
    .B2(_07087_),
    .X(_07335_));
 sky130_fd_sc_hd__nand4_1 _14646_ (.A(_07083_),
    .B(_07078_),
    .C(_07334_),
    .D(_07335_),
    .Y(_07336_));
 sky130_fd_sc_hd__a22o_1 _14647_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[5] ),
    .A2(_07078_),
    .B1(_07334_),
    .B2(_07335_),
    .X(_07337_));
 sky130_fd_sc_hd__nand2_1 _14648_ (.A(_07336_),
    .B(_07337_),
    .Y(_07338_));
 sky130_fd_sc_hd__and2_1 _14649_ (.A(_07291_),
    .B(_07294_),
    .X(_07339_));
 sky130_fd_sc_hd__xor2_2 _14650_ (.A(_07338_),
    .B(_07339_),
    .X(_07340_));
 sky130_fd_sc_hd__xor2_1 _14651_ (.A(_07332_),
    .B(_07340_),
    .X(_07341_));
 sky130_fd_sc_hd__o21ai_2 _14652_ (.A1(_07326_),
    .A2(_07327_),
    .B1(_07341_),
    .Y(_07342_));
 sky130_fd_sc_hd__or3_1 _14653_ (.A(_07326_),
    .B(_07327_),
    .C(_07341_),
    .X(_07343_));
 sky130_fd_sc_hd__nand3_1 _14654_ (.A(_07325_),
    .B(_07342_),
    .C(_07343_),
    .Y(_07344_));
 sky130_fd_sc_hd__a21o_1 _14655_ (.A1(_07342_),
    .A2(_07343_),
    .B1(_07325_),
    .X(_07345_));
 sky130_fd_sc_hd__and2_2 _14656_ (.A(_07344_),
    .B(_07345_),
    .X(_07346_));
 sky130_fd_sc_hd__nand2_1 _14657_ (.A(_07284_),
    .B(_07301_),
    .Y(_07347_));
 sky130_fd_sc_hd__o21ai_4 _14658_ (.A1(_07299_),
    .A2(_07300_),
    .B1(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__xnor2_4 _14659_ (.A(_07346_),
    .B(_07348_),
    .Y(_07349_));
 sky130_fd_sc_hd__xnor2_4 _14660_ (.A(_07318_),
    .B(_07349_),
    .Y(_07350_));
 sky130_fd_sc_hd__or2b_1 _14661_ (.A(_07302_),
    .B_N(_07303_),
    .X(_07351_));
 sky130_fd_sc_hd__or2b_1 _14662_ (.A(_07304_),
    .B_N(_07275_),
    .X(_07352_));
 sky130_fd_sc_hd__nand2_2 _14663_ (.A(_07351_),
    .B(_07352_),
    .Y(_07353_));
 sky130_fd_sc_hd__xor2_4 _14664_ (.A(_07350_),
    .B(_07353_),
    .X(_07354_));
 sky130_fd_sc_hd__xnor2_1 _14665_ (.A(_07316_),
    .B(_07354_),
    .Y(_07355_));
 sky130_fd_sc_hd__nor2_1 _14666_ (.A(_07314_),
    .B(_07355_),
    .Y(_07356_));
 sky130_fd_sc_hd__a21o_1 _14667_ (.A1(_07314_),
    .A2(_07355_),
    .B1(_07057_),
    .X(_07357_));
 sky130_fd_sc_hd__o221a_1 _14668_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[9] ),
    .A2(_07048_),
    .B1(_07356_),
    .B2(_07357_),
    .C1(_06180_),
    .X(_00432_));
 sky130_fd_sc_hd__a21o_1 _14669_ (.A1(_07308_),
    .A2(_07309_),
    .B1(_07354_),
    .X(_07358_));
 sky130_fd_sc_hd__a22oi_4 _14670_ (.A1(_07316_),
    .A2(_07354_),
    .B1(_07358_),
    .B2(_07314_),
    .Y(_07359_));
 sky130_fd_sc_hd__nand2_1 _14671_ (.A(_07350_),
    .B(_07353_),
    .Y(_07360_));
 sky130_fd_sc_hd__nand2_1 _14672_ (.A(_07346_),
    .B(_07348_),
    .Y(_07361_));
 sky130_fd_sc_hd__or2b_4 _14673_ (.A(_07349_),
    .B_N(_07318_),
    .X(_07362_));
 sky130_fd_sc_hd__o21bai_2 _14674_ (.A1(_07319_),
    .A2(_07323_),
    .B1_N(_07322_),
    .Y(_07363_));
 sky130_fd_sc_hd__clkbuf_4 _14675_ (.A(_07281_),
    .X(_07364_));
 sky130_fd_sc_hd__a21o_1 _14676_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[9] ),
    .A2(_07364_),
    .B1(_07280_),
    .X(_07365_));
 sky130_fd_sc_hd__xnor2_1 _14677_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[10] ),
    .B(_07281_),
    .Y(_07366_));
 sky130_fd_sc_hd__o21ai_1 _14678_ (.A1(_07328_),
    .A2(_07331_),
    .B1(_07330_),
    .Y(_07367_));
 sky130_fd_sc_hd__and2b_1 _14679_ (.A_N(_07366_),
    .B(_07367_),
    .X(_07368_));
 sky130_fd_sc_hd__and2b_1 _14680_ (.A_N(_07367_),
    .B(_07366_),
    .X(_07369_));
 sky130_fd_sc_hd__nor2_1 _14681_ (.A(_07368_),
    .B(_07369_),
    .Y(_07370_));
 sky130_fd_sc_hd__xor2_1 _14682_ (.A(_07365_),
    .B(_07370_),
    .X(_07371_));
 sky130_fd_sc_hd__or2_1 _14683_ (.A(_07338_),
    .B(_07339_),
    .X(_07372_));
 sky130_fd_sc_hd__nand2_1 _14684_ (.A(_07332_),
    .B(_07340_),
    .Y(_07373_));
 sky130_fd_sc_hd__a22o_1 _14685_ (.A1(_07079_),
    .A2(_07086_),
    .B1(_07090_),
    .B2(_07074_),
    .X(_07374_));
 sky130_fd_sc_hd__nand4_1 _14686_ (.A(_07079_),
    .B(_07074_),
    .C(_07086_),
    .D(_07090_),
    .Y(_07375_));
 sky130_fd_sc_hd__nand2_1 _14687_ (.A(_07374_),
    .B(_07375_),
    .Y(_07376_));
 sky130_fd_sc_hd__xor2_1 _14688_ (.A(_07328_),
    .B(_07376_),
    .X(_07377_));
 sky130_fd_sc_hd__inv_2 _14689_ (.A(_07078_),
    .Y(_07378_));
 sky130_fd_sc_hd__or4_1 _14690_ (.A(_07241_),
    .B(_07242_),
    .C(_07073_),
    .D(_07378_),
    .X(_07379_));
 sky130_fd_sc_hd__a22o_1 _14691_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[7] ),
    .A2(_07333_),
    .B1(_07078_),
    .B2(_07087_),
    .X(_07380_));
 sky130_fd_sc_hd__nand4_1 _14692_ (.A(_07083_),
    .B(_07082_),
    .C(_07379_),
    .D(_07380_),
    .Y(_07381_));
 sky130_fd_sc_hd__a22o_1 _14693_ (.A1(_07083_),
    .A2(_07082_),
    .B1(_07379_),
    .B2(_07380_),
    .X(_07382_));
 sky130_fd_sc_hd__nand2_1 _14694_ (.A(_07381_),
    .B(_07382_),
    .Y(_07383_));
 sky130_fd_sc_hd__nand2_1 _14695_ (.A(_07334_),
    .B(_07336_),
    .Y(_07384_));
 sky130_fd_sc_hd__xnor2_1 _14696_ (.A(_07383_),
    .B(_07384_),
    .Y(_07385_));
 sky130_fd_sc_hd__xnor2_1 _14697_ (.A(_07377_),
    .B(_07385_),
    .Y(_07386_));
 sky130_fd_sc_hd__a21o_1 _14698_ (.A1(_07372_),
    .A2(_07373_),
    .B1(_07386_),
    .X(_07387_));
 sky130_fd_sc_hd__nand3_1 _14699_ (.A(_07372_),
    .B(_07373_),
    .C(_07386_),
    .Y(_07388_));
 sky130_fd_sc_hd__nand3_1 _14700_ (.A(_07371_),
    .B(_07387_),
    .C(_07388_),
    .Y(_07389_));
 sky130_fd_sc_hd__inv_2 _14701_ (.A(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__a21oi_1 _14702_ (.A1(_07387_),
    .A2(_07388_),
    .B1(_07371_),
    .Y(_07391_));
 sky130_fd_sc_hd__a211o_1 _14703_ (.A1(_07342_),
    .A2(_07344_),
    .B1(_07390_),
    .C1(_07391_),
    .X(_07392_));
 sky130_fd_sc_hd__o211ai_2 _14704_ (.A1(_07390_),
    .A2(_07391_),
    .B1(_07342_),
    .C1(_07344_),
    .Y(_07393_));
 sky130_fd_sc_hd__and3_1 _14705_ (.A(_07363_),
    .B(_07392_),
    .C(_07393_),
    .X(_07394_));
 sky130_fd_sc_hd__a21oi_2 _14706_ (.A1(_07392_),
    .A2(_07393_),
    .B1(_07363_),
    .Y(_07395_));
 sky130_fd_sc_hd__a211oi_2 _14707_ (.A1(_07361_),
    .A2(_07362_),
    .B1(_07394_),
    .C1(_07395_),
    .Y(_07396_));
 sky130_fd_sc_hd__o211a_1 _14708_ (.A1(_07394_),
    .A2(_07395_),
    .B1(_07361_),
    .C1(_07362_),
    .X(_07397_));
 sky130_fd_sc_hd__or3_4 _14709_ (.A(_07360_),
    .B(_07396_),
    .C(_07397_),
    .X(_07398_));
 sky130_fd_sc_hd__o21ai_1 _14710_ (.A1(_07396_),
    .A2(_07397_),
    .B1(_07360_),
    .Y(_07399_));
 sky130_fd_sc_hd__and2_1 _14711_ (.A(_07398_),
    .B(_07399_),
    .X(_07400_));
 sky130_fd_sc_hd__xnor2_1 _14712_ (.A(_07359_),
    .B(_07400_),
    .Y(_07401_));
 sky130_fd_sc_hd__or2_1 _14713_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[10] ),
    .B(_06168_),
    .X(_07402_));
 sky130_fd_sc_hd__o211a_1 _14714_ (.A1(_06848_),
    .A2(_07401_),
    .B1(_07402_),
    .C1(_07092_),
    .X(_00433_));
 sky130_fd_sc_hd__or2b_1 _14715_ (.A(_07359_),
    .B_N(_07400_),
    .X(_07403_));
 sky130_fd_sc_hd__a21o_1 _14716_ (.A1(_07365_),
    .A2(_07370_),
    .B1(_07368_),
    .X(_07404_));
 sky130_fd_sc_hd__a21o_1 _14717_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[10] ),
    .A2(_07364_),
    .B1(_07280_),
    .X(_07405_));
 sky130_fd_sc_hd__o21ai_1 _14718_ (.A1(_07328_),
    .A2(_07376_),
    .B1(_07375_),
    .Y(_07406_));
 sky130_fd_sc_hd__xnor2_1 _14719_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[11] ),
    .B(_07281_),
    .Y(_07407_));
 sky130_fd_sc_hd__xnor2_1 _14720_ (.A(_07406_),
    .B(_07407_),
    .Y(_07408_));
 sky130_fd_sc_hd__xnor2_1 _14721_ (.A(_07405_),
    .B(_07408_),
    .Y(_07409_));
 sky130_fd_sc_hd__or2b_1 _14722_ (.A(_07383_),
    .B_N(_07384_),
    .X(_07410_));
 sky130_fd_sc_hd__nand2_1 _14723_ (.A(_07377_),
    .B(_07385_),
    .Y(_07411_));
 sky130_fd_sc_hd__and3_1 _14724_ (.A(_07079_),
    .B(_07074_),
    .C(_07089_),
    .X(_07412_));
 sky130_fd_sc_hd__o21ai_1 _14725_ (.A1(_07079_),
    .A2(_07074_),
    .B1(_07090_),
    .Y(_07413_));
 sky130_fd_sc_hd__nor2_2 _14726_ (.A(_07412_),
    .B(_07413_),
    .Y(_07414_));
 sky130_fd_sc_hd__xnor2_4 _14727_ (.A(_07328_),
    .B(_07414_),
    .Y(_07415_));
 sky130_fd_sc_hd__inv_2 _14728_ (.A(net1123),
    .Y(_07416_));
 sky130_fd_sc_hd__or4_1 _14729_ (.A(_07241_),
    .B(_07242_),
    .C(_07078_),
    .D(_07416_),
    .X(_07417_));
 sky130_fd_sc_hd__a22o_1 _14730_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[7] ),
    .A2(_07378_),
    .B1(_07082_),
    .B2(_07087_),
    .X(_07418_));
 sky130_fd_sc_hd__nand4_1 _14731_ (.A(_07083_),
    .B(_07086_),
    .C(_07417_),
    .D(_07418_),
    .Y(_07419_));
 sky130_fd_sc_hd__a22o_1 _14732_ (.A1(_07083_),
    .A2(_07086_),
    .B1(_07417_),
    .B2(_07418_),
    .X(_07420_));
 sky130_fd_sc_hd__nand2_1 _14733_ (.A(_07419_),
    .B(_07420_),
    .Y(_07421_));
 sky130_fd_sc_hd__nand2_1 _14734_ (.A(_07379_),
    .B(_07381_),
    .Y(_07422_));
 sky130_fd_sc_hd__xnor2_1 _14735_ (.A(_07421_),
    .B(_07422_),
    .Y(_07423_));
 sky130_fd_sc_hd__xnor2_1 _14736_ (.A(_07415_),
    .B(_07423_),
    .Y(_07424_));
 sky130_fd_sc_hd__a21o_1 _14737_ (.A1(_07410_),
    .A2(_07411_),
    .B1(_07424_),
    .X(_07425_));
 sky130_fd_sc_hd__nand3_1 _14738_ (.A(_07410_),
    .B(_07411_),
    .C(_07424_),
    .Y(_07426_));
 sky130_fd_sc_hd__nand2_1 _14739_ (.A(_07425_),
    .B(_07426_),
    .Y(_07427_));
 sky130_fd_sc_hd__or2_1 _14740_ (.A(_07409_),
    .B(_07427_),
    .X(_07428_));
 sky130_fd_sc_hd__nand2_1 _14741_ (.A(_07409_),
    .B(_07427_),
    .Y(_07429_));
 sky130_fd_sc_hd__nand2_1 _14742_ (.A(_07387_),
    .B(_07389_),
    .Y(_07430_));
 sky130_fd_sc_hd__nand3_1 _14743_ (.A(_07428_),
    .B(_07429_),
    .C(_07430_),
    .Y(_07431_));
 sky130_fd_sc_hd__a21o_1 _14744_ (.A1(_07428_),
    .A2(_07429_),
    .B1(_07430_),
    .X(_07432_));
 sky130_fd_sc_hd__nand2_1 _14745_ (.A(_07431_),
    .B(_07432_),
    .Y(_07433_));
 sky130_fd_sc_hd__xor2_1 _14746_ (.A(_07404_),
    .B(_07433_),
    .X(_07434_));
 sky130_fd_sc_hd__a21bo_1 _14747_ (.A1(_07363_),
    .A2(_07393_),
    .B1_N(_07392_),
    .X(_07435_));
 sky130_fd_sc_hd__xor2_1 _14748_ (.A(_07434_),
    .B(_07435_),
    .X(_07436_));
 sky130_fd_sc_hd__xnor2_1 _14749_ (.A(_07396_),
    .B(_07436_),
    .Y(_07437_));
 sky130_fd_sc_hd__a21oi_1 _14750_ (.A1(_07398_),
    .A2(_07403_),
    .B1(net1124),
    .Y(_07438_));
 sky130_fd_sc_hd__clkbuf_8 _14751_ (.A(_05633_),
    .X(_07439_));
 sky130_fd_sc_hd__a31o_1 _14752_ (.A1(_07398_),
    .A2(_07403_),
    .A3(net1124),
    .B1(_07439_),
    .X(_07440_));
 sky130_fd_sc_hd__o221a_1 _14753_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[11] ),
    .A2(_07048_),
    .B1(_07438_),
    .B2(_07440_),
    .C1(_06180_),
    .X(_00434_));
 sky130_fd_sc_hd__and2b_1 _14754_ (.A_N(_07437_),
    .B(_07359_),
    .X(_07441_));
 sky130_fd_sc_hd__a211o_1 _14755_ (.A1(_07361_),
    .A2(_07362_),
    .B1(_07394_),
    .C1(_07395_),
    .X(_07442_));
 sky130_fd_sc_hd__a21oi_1 _14756_ (.A1(_07442_),
    .A2(_07398_),
    .B1(_07436_),
    .Y(_07443_));
 sky130_fd_sc_hd__a21o_1 _14757_ (.A1(_07400_),
    .A2(_07441_),
    .B1(_07443_),
    .X(_07444_));
 sky130_fd_sc_hd__or2b_1 _14758_ (.A(_07434_),
    .B_N(_07435_),
    .X(_07445_));
 sky130_fd_sc_hd__a21bo_1 _14759_ (.A1(_07404_),
    .A2(_07432_),
    .B1_N(_07431_),
    .X(_07446_));
 sky130_fd_sc_hd__or2b_1 _14760_ (.A(_07407_),
    .B_N(_07406_),
    .X(_07447_));
 sky130_fd_sc_hd__a21bo_1 _14761_ (.A1(_07405_),
    .A2(_07408_),
    .B1_N(_07447_),
    .X(_07448_));
 sky130_fd_sc_hd__a21o_1 _14762_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[11] ),
    .A2(_07364_),
    .B1(_07280_),
    .X(_07449_));
 sky130_fd_sc_hd__o21ba_2 _14763_ (.A1(_07328_),
    .A2(_07413_),
    .B1_N(_07412_),
    .X(_07450_));
 sky130_fd_sc_hd__xnor2_1 _14764_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[12] ),
    .B(_07281_),
    .Y(_07451_));
 sky130_fd_sc_hd__nor2_1 _14765_ (.A(_07450_),
    .B(_07451_),
    .Y(_07452_));
 sky130_fd_sc_hd__and2_1 _14766_ (.A(_07450_),
    .B(_07451_),
    .X(_07453_));
 sky130_fd_sc_hd__nor2_1 _14767_ (.A(_07452_),
    .B(_07453_),
    .Y(_07454_));
 sky130_fd_sc_hd__xnor2_1 _14768_ (.A(_07449_),
    .B(_07454_),
    .Y(_07455_));
 sky130_fd_sc_hd__or2b_1 _14769_ (.A(_07421_),
    .B_N(_07422_),
    .X(_07456_));
 sky130_fd_sc_hd__nand2_1 _14770_ (.A(_07415_),
    .B(_07423_),
    .Y(_07457_));
 sky130_fd_sc_hd__nand2_1 _14771_ (.A(_07417_),
    .B(_07419_),
    .Y(_07458_));
 sky130_fd_sc_hd__nand2_2 _14772_ (.A(_07083_),
    .B(_07090_),
    .Y(_07459_));
 sky130_fd_sc_hd__inv_2 _14773_ (.A(_07085_),
    .Y(_07460_));
 sky130_fd_sc_hd__or4_4 _14774_ (.A(_07241_),
    .B(_07242_),
    .C(_07082_),
    .D(_07460_),
    .X(_07461_));
 sky130_fd_sc_hd__a22o_1 _14775_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[7] ),
    .A2(_07416_),
    .B1(_07085_),
    .B2(_07087_),
    .X(_07462_));
 sky130_fd_sc_hd__nand2_2 _14776_ (.A(_07461_),
    .B(_07462_),
    .Y(_07463_));
 sky130_fd_sc_hd__xnor2_1 _14777_ (.A(_07459_),
    .B(_07463_),
    .Y(_07464_));
 sky130_fd_sc_hd__xnor2_1 _14778_ (.A(_07458_),
    .B(_07464_),
    .Y(_07465_));
 sky130_fd_sc_hd__xnor2_1 _14779_ (.A(_07415_),
    .B(_07465_),
    .Y(_07466_));
 sky130_fd_sc_hd__a21o_1 _14780_ (.A1(_07456_),
    .A2(_07457_),
    .B1(_07466_),
    .X(_07467_));
 sky130_fd_sc_hd__nand3_1 _14781_ (.A(_07456_),
    .B(_07457_),
    .C(_07466_),
    .Y(_07468_));
 sky130_fd_sc_hd__nand2_1 _14782_ (.A(_07467_),
    .B(_07468_),
    .Y(_07469_));
 sky130_fd_sc_hd__or2_1 _14783_ (.A(_07455_),
    .B(_07469_),
    .X(_07470_));
 sky130_fd_sc_hd__inv_2 _14784_ (.A(_07470_),
    .Y(_07471_));
 sky130_fd_sc_hd__and2_1 _14785_ (.A(_07455_),
    .B(_07469_),
    .X(_07472_));
 sky130_fd_sc_hd__a211o_1 _14786_ (.A1(_07425_),
    .A2(_07428_),
    .B1(_07471_),
    .C1(_07472_),
    .X(_07473_));
 sky130_fd_sc_hd__o211ai_1 _14787_ (.A1(_07471_),
    .A2(_07472_),
    .B1(_07425_),
    .C1(_07428_),
    .Y(_07474_));
 sky130_fd_sc_hd__and3_1 _14788_ (.A(_07448_),
    .B(_07473_),
    .C(_07474_),
    .X(_07475_));
 sky130_fd_sc_hd__a21oi_1 _14789_ (.A1(_07473_),
    .A2(_07474_),
    .B1(_07448_),
    .Y(_07476_));
 sky130_fd_sc_hd__or2_1 _14790_ (.A(_07475_),
    .B(_07476_),
    .X(_07477_));
 sky130_fd_sc_hd__xnor2_2 _14791_ (.A(_07446_),
    .B(_07477_),
    .Y(_07478_));
 sky130_fd_sc_hd__xnor2_1 _14792_ (.A(_07445_),
    .B(_07478_),
    .Y(_07479_));
 sky130_fd_sc_hd__nand2_1 _14793_ (.A(_07444_),
    .B(_07479_),
    .Y(_07480_));
 sky130_fd_sc_hd__or2_1 _14794_ (.A(_07444_),
    .B(_07479_),
    .X(_07481_));
 sky130_fd_sc_hd__a21o_1 _14795_ (.A1(_07480_),
    .A2(_07481_),
    .B1(_06682_),
    .X(_07482_));
 sky130_fd_sc_hd__o211a_1 _14796_ (.A1(net1065),
    .A2(_06660_),
    .B1(_07482_),
    .C1(_07092_),
    .X(_00435_));
 sky130_fd_sc_hd__or2b_4 _14797_ (.A(_07445_),
    .B_N(_07478_),
    .X(_07483_));
 sky130_fd_sc_hd__or2b_4 _14798_ (.A(_07477_),
    .B_N(_07446_),
    .X(_07484_));
 sky130_fd_sc_hd__inv_2 _14799_ (.A(_07473_),
    .Y(_07485_));
 sky130_fd_sc_hd__a21o_1 _14800_ (.A1(_07449_),
    .A2(_07454_),
    .B1(_07452_),
    .X(_07486_));
 sky130_fd_sc_hd__a21o_1 _14801_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[12] ),
    .A2(_07364_),
    .B1(_07280_),
    .X(_07487_));
 sky130_fd_sc_hd__xnor2_1 _14802_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[13] ),
    .B(_07364_),
    .Y(_07488_));
 sky130_fd_sc_hd__nor2_1 _14803_ (.A(_07450_),
    .B(_07488_),
    .Y(_07489_));
 sky130_fd_sc_hd__and2_1 _14804_ (.A(_07450_),
    .B(_07488_),
    .X(_07490_));
 sky130_fd_sc_hd__nor2_1 _14805_ (.A(_07489_),
    .B(_07490_),
    .Y(_07491_));
 sky130_fd_sc_hd__xnor2_1 _14806_ (.A(_07487_),
    .B(_07491_),
    .Y(_07492_));
 sky130_fd_sc_hd__or2b_1 _14807_ (.A(_07464_),
    .B_N(_07458_),
    .X(_07493_));
 sky130_fd_sc_hd__nand2_1 _14808_ (.A(_07415_),
    .B(_07465_),
    .Y(_07494_));
 sky130_fd_sc_hd__o21ai_1 _14809_ (.A1(_07459_),
    .A2(_07463_),
    .B1(_07461_),
    .Y(_07495_));
 sky130_fd_sc_hd__nand2_1 _14810_ (.A(_07087_),
    .B(_07089_),
    .Y(_07496_));
 sky130_fd_sc_hd__or3_1 _14811_ (.A(_07241_),
    .B(_07085_),
    .C(_07496_),
    .X(_07497_));
 sky130_fd_sc_hd__o21ai_1 _14812_ (.A1(_07241_),
    .A2(_07086_),
    .B1(_07496_),
    .Y(_07498_));
 sky130_fd_sc_hd__nand2_1 _14813_ (.A(_07497_),
    .B(_07498_),
    .Y(_07499_));
 sky130_fd_sc_hd__xnor2_1 _14814_ (.A(_07459_),
    .B(_07499_),
    .Y(_07500_));
 sky130_fd_sc_hd__xnor2_1 _14815_ (.A(_07495_),
    .B(_07500_),
    .Y(_07501_));
 sky130_fd_sc_hd__and2_1 _14816_ (.A(_07415_),
    .B(_07501_),
    .X(_07502_));
 sky130_fd_sc_hd__nor2_1 _14817_ (.A(_07415_),
    .B(_07501_),
    .Y(_07503_));
 sky130_fd_sc_hd__or2_1 _14818_ (.A(_07502_),
    .B(_07503_),
    .X(_07504_));
 sky130_fd_sc_hd__a21o_1 _14819_ (.A1(_07493_),
    .A2(_07494_),
    .B1(_07504_),
    .X(_07505_));
 sky130_fd_sc_hd__nand3_1 _14820_ (.A(_07493_),
    .B(_07494_),
    .C(_07504_),
    .Y(_07506_));
 sky130_fd_sc_hd__nand2_1 _14821_ (.A(_07505_),
    .B(_07506_),
    .Y(_07507_));
 sky130_fd_sc_hd__xnor2_1 _14822_ (.A(_07492_),
    .B(_07507_),
    .Y(_07508_));
 sky130_fd_sc_hd__a21o_1 _14823_ (.A1(_07467_),
    .A2(_07470_),
    .B1(_07508_),
    .X(_07509_));
 sky130_fd_sc_hd__nand3_1 _14824_ (.A(_07467_),
    .B(_07470_),
    .C(_07508_),
    .Y(_07510_));
 sky130_fd_sc_hd__and3_1 _14825_ (.A(_07486_),
    .B(_07509_),
    .C(_07510_),
    .X(_07511_));
 sky130_fd_sc_hd__a21oi_1 _14826_ (.A1(_07509_),
    .A2(_07510_),
    .B1(_07486_),
    .Y(_07512_));
 sky130_fd_sc_hd__nor2_1 _14827_ (.A(_07511_),
    .B(_07512_),
    .Y(_07513_));
 sky130_fd_sc_hd__o21ai_1 _14828_ (.A1(_07485_),
    .A2(_07475_),
    .B1(_07513_),
    .Y(_07514_));
 sky130_fd_sc_hd__or3_1 _14829_ (.A(_07485_),
    .B(_07475_),
    .C(_07513_),
    .X(_07515_));
 sky130_fd_sc_hd__nand2_1 _14830_ (.A(_07514_),
    .B(_07515_),
    .Y(_07516_));
 sky130_fd_sc_hd__xor2_2 _14831_ (.A(_07484_),
    .B(_07516_),
    .X(_07517_));
 sky130_fd_sc_hd__a21oi_1 _14832_ (.A1(_07483_),
    .A2(_07480_),
    .B1(_07517_),
    .Y(_07518_));
 sky130_fd_sc_hd__a31o_1 _14833_ (.A1(_07483_),
    .A2(_07480_),
    .A3(_07517_),
    .B1(_07439_),
    .X(_07519_));
 sky130_fd_sc_hd__o221a_1 _14834_ (.A1(net1066),
    .A2(_07048_),
    .B1(_07518_),
    .B2(_07519_),
    .C1(_06180_),
    .X(_00436_));
 sky130_fd_sc_hd__a21bo_1 _14835_ (.A1(_07486_),
    .A2(_07510_),
    .B1_N(_07509_),
    .X(_07520_));
 sky130_fd_sc_hd__a21o_1 _14836_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[13] ),
    .A2(_07364_),
    .B1(_07280_),
    .X(_07521_));
 sky130_fd_sc_hd__xnor2_1 _14837_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[14] ),
    .B(_07364_),
    .Y(_07522_));
 sky130_fd_sc_hd__nor2_1 _14838_ (.A(_07450_),
    .B(_07522_),
    .Y(_07523_));
 sky130_fd_sc_hd__and2_1 _14839_ (.A(_07450_),
    .B(_07522_),
    .X(_07524_));
 sky130_fd_sc_hd__nor2_1 _14840_ (.A(_07523_),
    .B(_07524_),
    .Y(_07525_));
 sky130_fd_sc_hd__xnor2_1 _14841_ (.A(_07521_),
    .B(_07525_),
    .Y(_07526_));
 sky130_fd_sc_hd__and2b_1 _14842_ (.A_N(_07500_),
    .B(_07495_),
    .X(_07527_));
 sky130_fd_sc_hd__o211a_1 _14843_ (.A1(_07241_),
    .A2(_07090_),
    .B1(_07459_),
    .C1(_07496_),
    .X(_07528_));
 sky130_fd_sc_hd__o21a_1 _14844_ (.A1(_07459_),
    .A2(_07499_),
    .B1(_07497_),
    .X(_07529_));
 sky130_fd_sc_hd__a31oi_2 _14845_ (.A1(_07087_),
    .A2(_07083_),
    .A3(_07090_),
    .B1(_07529_),
    .Y(_07530_));
 sky130_fd_sc_hd__inv_2 _14846_ (.A(_07415_),
    .Y(_07531_));
 sky130_fd_sc_hd__o21a_1 _14847_ (.A1(_07528_),
    .A2(_07530_),
    .B1(_07531_),
    .X(_07532_));
 sky130_fd_sc_hd__or3_1 _14848_ (.A(_07531_),
    .B(_07528_),
    .C(_07530_),
    .X(_07533_));
 sky130_fd_sc_hd__or2b_1 _14849_ (.A(_07532_),
    .B_N(_07533_),
    .X(_07534_));
 sky130_fd_sc_hd__o21ba_1 _14850_ (.A1(_07527_),
    .A2(_07502_),
    .B1_N(_07534_),
    .X(_07535_));
 sky130_fd_sc_hd__or3b_1 _14851_ (.A(_07527_),
    .B(_07502_),
    .C_N(_07534_),
    .X(_07536_));
 sky130_fd_sc_hd__and2b_1 _14852_ (.A_N(_07535_),
    .B(_07536_),
    .X(_07537_));
 sky130_fd_sc_hd__xor2_1 _14853_ (.A(_07526_),
    .B(_07537_),
    .X(_07538_));
 sky130_fd_sc_hd__o21a_1 _14854_ (.A1(_07492_),
    .A2(_07507_),
    .B1(_07505_),
    .X(_07539_));
 sky130_fd_sc_hd__or2_1 _14855_ (.A(_07538_),
    .B(_07539_),
    .X(_07540_));
 sky130_fd_sc_hd__nand2_1 _14856_ (.A(_07538_),
    .B(_07539_),
    .Y(_07541_));
 sky130_fd_sc_hd__nand2_1 _14857_ (.A(_07540_),
    .B(_07541_),
    .Y(_07542_));
 sky130_fd_sc_hd__a21o_1 _14858_ (.A1(_07487_),
    .A2(_07491_),
    .B1(_07489_),
    .X(_07543_));
 sky130_fd_sc_hd__or2b_1 _14859_ (.A(_07542_),
    .B_N(_07543_),
    .X(_07544_));
 sky130_fd_sc_hd__or2b_1 _14860_ (.A(_07543_),
    .B_N(_07542_),
    .X(_07545_));
 sky130_fd_sc_hd__nand2_1 _14861_ (.A(_07544_),
    .B(_07545_),
    .Y(_07546_));
 sky130_fd_sc_hd__xor2_1 _14862_ (.A(_07520_),
    .B(_07546_),
    .X(_07547_));
 sky130_fd_sc_hd__or2_1 _14863_ (.A(_07514_),
    .B(_07547_),
    .X(_07548_));
 sky130_fd_sc_hd__nand2_1 _14864_ (.A(_07514_),
    .B(_07547_),
    .Y(_07549_));
 sky130_fd_sc_hd__and2_1 _14865_ (.A(_07548_),
    .B(_07549_),
    .X(_07550_));
 sky130_fd_sc_hd__a21oi_1 _14866_ (.A1(_07484_),
    .A2(_07483_),
    .B1(_07516_),
    .Y(_07551_));
 sky130_fd_sc_hd__a31o_1 _14867_ (.A1(_07444_),
    .A2(_07479_),
    .A3(_07517_),
    .B1(_07551_),
    .X(_07552_));
 sky130_fd_sc_hd__nand2_1 _14868_ (.A(_07550_),
    .B(_07552_),
    .Y(_07553_));
 sky130_fd_sc_hd__or2_1 _14869_ (.A(_07550_),
    .B(_07552_),
    .X(_07554_));
 sky130_fd_sc_hd__a21o_1 _14870_ (.A1(_07553_),
    .A2(_07554_),
    .B1(_06682_),
    .X(_07555_));
 sky130_fd_sc_hd__o211a_1 _14871_ (.A1(net1062),
    .A2(_06660_),
    .B1(_07555_),
    .C1(_07092_),
    .X(_00437_));
 sky130_fd_sc_hd__inv_2 _14872_ (.A(_07548_),
    .Y(_07556_));
 sky130_fd_sc_hd__a21oi_1 _14873_ (.A1(_07550_),
    .A2(_07552_),
    .B1(_07556_),
    .Y(_07557_));
 sky130_fd_sc_hd__and2b_1 _14874_ (.A_N(_07546_),
    .B(_07520_),
    .X(_07558_));
 sky130_fd_sc_hd__a21o_1 _14875_ (.A1(_07521_),
    .A2(_07525_),
    .B1(_07523_),
    .X(_07559_));
 sky130_fd_sc_hd__and2b_1 _14876_ (.A_N(_07526_),
    .B(_07537_),
    .X(_07560_));
 sky130_fd_sc_hd__a21oi_1 _14877_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[14] ),
    .A2(_07364_),
    .B1(_07280_),
    .Y(_07561_));
 sky130_fd_sc_hd__xnor2_2 _14878_ (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[15] ),
    .B(_07364_),
    .Y(_07562_));
 sky130_fd_sc_hd__xor2_2 _14879_ (.A(_07450_),
    .B(_07562_),
    .X(_07563_));
 sky130_fd_sc_hd__xor2_1 _14880_ (.A(_07561_),
    .B(_07563_),
    .X(_07564_));
 sky130_fd_sc_hd__xor2_1 _14881_ (.A(_07532_),
    .B(_07564_),
    .X(_07565_));
 sky130_fd_sc_hd__o21a_1 _14882_ (.A1(_07535_),
    .A2(_07560_),
    .B1(_07565_),
    .X(_07566_));
 sky130_fd_sc_hd__nor3_1 _14883_ (.A(_07535_),
    .B(_07560_),
    .C(_07565_),
    .Y(_07567_));
 sky130_fd_sc_hd__nor2_1 _14884_ (.A(_07566_),
    .B(_07567_),
    .Y(_07568_));
 sky130_fd_sc_hd__xnor2_1 _14885_ (.A(_07559_),
    .B(_07568_),
    .Y(_07569_));
 sky130_fd_sc_hd__a21o_1 _14886_ (.A1(_07540_),
    .A2(_07544_),
    .B1(_07569_),
    .X(_07570_));
 sky130_fd_sc_hd__nand3_1 _14887_ (.A(_07540_),
    .B(_07544_),
    .C(_07569_),
    .Y(_07571_));
 sky130_fd_sc_hd__and2_1 _14888_ (.A(_07570_),
    .B(_07571_),
    .X(_07572_));
 sky130_fd_sc_hd__xor2_2 _14889_ (.A(_07558_),
    .B(_07572_),
    .X(_07573_));
 sky130_fd_sc_hd__nor2_1 _14890_ (.A(_07557_),
    .B(_07573_),
    .Y(_07574_));
 sky130_fd_sc_hd__a21o_1 _14891_ (.A1(_07557_),
    .A2(_07573_),
    .B1(_07057_),
    .X(_07575_));
 sky130_fd_sc_hd__o221a_1 _14892_ (.A1(net1088),
    .A2(_07048_),
    .B1(_07574_),
    .B2(_07575_),
    .C1(_06180_),
    .X(_00438_));
 sky130_fd_sc_hd__buf_8 _14893_ (.A(_05731_),
    .X(_07576_));
 sky130_fd_sc_hd__and2_1 _14894_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[16] ),
    .B(_07576_),
    .X(_07577_));
 sky130_fd_sc_hd__and3_1 _14895_ (.A(_07550_),
    .B(_07552_),
    .C(_07573_),
    .X(_07578_));
 sky130_fd_sc_hd__a21o_1 _14896_ (.A1(_07559_),
    .A2(_07568_),
    .B1(_07566_),
    .X(_07579_));
 sky130_fd_sc_hd__or2b_1 _14897_ (.A(_07561_),
    .B_N(_07563_),
    .X(_07580_));
 sky130_fd_sc_hd__o21ai_1 _14898_ (.A1(_07450_),
    .A2(_07562_),
    .B1(_07580_),
    .Y(_07581_));
 sky130_fd_sc_hd__and2_1 _14899_ (.A(_07531_),
    .B(_07528_),
    .X(_07582_));
 sky130_fd_sc_hd__a21oi_1 _14900_ (.A1(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[15] ),
    .A2(_07364_),
    .B1(_07280_),
    .Y(_07583_));
 sky130_fd_sc_hd__xnor2_1 _14901_ (.A(_07563_),
    .B(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__xnor2_1 _14902_ (.A(_07582_),
    .B(_07584_),
    .Y(_07585_));
 sky130_fd_sc_hd__o2bb2a_1 _14903_ (.A1_N(_07531_),
    .A2_N(_07530_),
    .B1(_07564_),
    .B2(_07582_),
    .X(_07586_));
 sky130_fd_sc_hd__xnor2_1 _14904_ (.A(_07585_),
    .B(_07586_),
    .Y(_07587_));
 sky130_fd_sc_hd__xnor2_1 _14905_ (.A(_07581_),
    .B(_07587_),
    .Y(_07588_));
 sky130_fd_sc_hd__xnor2_1 _14906_ (.A(_07579_),
    .B(_07588_),
    .Y(_07589_));
 sky130_fd_sc_hd__xnor2_1 _14907_ (.A(_07570_),
    .B(_07589_),
    .Y(_07590_));
 sky130_fd_sc_hd__o21ai_1 _14908_ (.A1(_07558_),
    .A2(_07556_),
    .B1(_07572_),
    .Y(_07591_));
 sky130_fd_sc_hd__and4b_2 _14909_ (.A_N(_07578_),
    .B(_07590_),
    .C(_07591_),
    .D(_05315_),
    .X(_07592_));
 sky130_fd_sc_hd__buf_6 _14910_ (.A(_07592_),
    .X(_07593_));
 sky130_fd_sc_hd__buf_2 _14911_ (.A(_05352_),
    .X(_07594_));
 sky130_fd_sc_hd__o21a_1 _14912_ (.A1(_07577_),
    .A2(net229),
    .B1(_07594_),
    .X(_00439_));
 sky130_fd_sc_hd__buf_8 _14913_ (.A(_05633_),
    .X(_07595_));
 sky130_fd_sc_hd__and2_1 _14914_ (.A(net1082),
    .B(_07595_),
    .X(_07596_));
 sky130_fd_sc_hd__o21a_1 _14915_ (.A1(net229),
    .A2(_07596_),
    .B1(_07594_),
    .X(_00440_));
 sky130_fd_sc_hd__and2_1 _14916_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[18] ),
    .B(_07595_),
    .X(_07597_));
 sky130_fd_sc_hd__o21a_1 _14917_ (.A1(net229),
    .A2(_07597_),
    .B1(_07594_),
    .X(_00441_));
 sky130_fd_sc_hd__and2_1 _14918_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[19] ),
    .B(_07595_),
    .X(_07598_));
 sky130_fd_sc_hd__o21a_1 _14919_ (.A1(net229),
    .A2(_07598_),
    .B1(_07594_),
    .X(_00442_));
 sky130_fd_sc_hd__and2_1 _14920_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[20] ),
    .B(_07595_),
    .X(_07599_));
 sky130_fd_sc_hd__o21a_1 _14921_ (.A1(net229),
    .A2(_07599_),
    .B1(_07594_),
    .X(_00443_));
 sky130_fd_sc_hd__and2_1 _14922_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[21] ),
    .B(_07595_),
    .X(_07600_));
 sky130_fd_sc_hd__o21a_1 _14923_ (.A1(_07593_),
    .A2(_07600_),
    .B1(_07594_),
    .X(_00444_));
 sky130_fd_sc_hd__and2_1 _14924_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[23] ),
    .B(_07595_),
    .X(_07601_));
 sky130_fd_sc_hd__o21a_1 _14925_ (.A1(_07593_),
    .A2(_07601_),
    .B1(_07594_),
    .X(_00445_));
 sky130_fd_sc_hd__and2_1 _14926_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[24] ),
    .B(_07576_),
    .X(_07602_));
 sky130_fd_sc_hd__o21a_1 _14927_ (.A1(_07593_),
    .A2(_07602_),
    .B1(_07594_),
    .X(_00446_));
 sky130_fd_sc_hd__and2_1 _14928_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[25] ),
    .B(_07576_),
    .X(_07603_));
 sky130_fd_sc_hd__o21a_1 _14929_ (.A1(_07593_),
    .A2(_07603_),
    .B1(_07594_),
    .X(_00447_));
 sky130_fd_sc_hd__and2_1 _14930_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[27] ),
    .B(_07576_),
    .X(_07604_));
 sky130_fd_sc_hd__o21a_1 _14931_ (.A1(_07593_),
    .A2(_07604_),
    .B1(_07594_),
    .X(_00448_));
 sky130_fd_sc_hd__and2_1 _14932_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[31] ),
    .B(_07576_),
    .X(_07605_));
 sky130_fd_sc_hd__o21a_1 _14933_ (.A1(_07592_),
    .A2(_07605_),
    .B1(_04870_),
    .X(_00449_));
 sky130_fd_sc_hd__clkbuf_4 _14934_ (.A(\top_inst.grid_inst.data_path_wires[6][0] ),
    .X(_07606_));
 sky130_fd_sc_hd__or2_1 _14935_ (.A(_05736_),
    .B(_07061_),
    .X(_07607_));
 sky130_fd_sc_hd__o211a_1 _14936_ (.A1(_07606_),
    .A2(_05735_),
    .B1(_07607_),
    .C1(_07092_),
    .X(_00450_));
 sky130_fd_sc_hd__clkbuf_4 _14937_ (.A(\top_inst.grid_inst.data_path_wires[6][1] ),
    .X(_07608_));
 sky130_fd_sc_hd__nand2_1 _14938_ (.A(_05739_),
    .B(_07292_),
    .Y(_07609_));
 sky130_fd_sc_hd__o211a_1 _14939_ (.A1(_07608_),
    .A2(_05735_),
    .B1(_07609_),
    .C1(_07092_),
    .X(_00451_));
 sky130_fd_sc_hd__clkbuf_4 _14940_ (.A(\top_inst.grid_inst.data_path_wires[6][2] ),
    .X(_07610_));
 sky130_fd_sc_hd__clkbuf_4 _14941_ (.A(_04865_),
    .X(_07611_));
 sky130_fd_sc_hd__nand2_1 _14942_ (.A(_05739_),
    .B(_07290_),
    .Y(_07612_));
 sky130_fd_sc_hd__o211a_1 _14943_ (.A1(_07610_),
    .A2(_07611_),
    .B1(_07612_),
    .C1(_07092_),
    .X(_00452_));
 sky130_fd_sc_hd__clkbuf_4 _14944_ (.A(\top_inst.grid_inst.data_path_wires[6][3] ),
    .X(_07613_));
 sky130_fd_sc_hd__nand2_1 _14945_ (.A(_04865_),
    .B(_07333_),
    .Y(_07614_));
 sky130_fd_sc_hd__o211a_1 _14946_ (.A1(_07613_),
    .A2(_07611_),
    .B1(_07614_),
    .C1(_07092_),
    .X(_00453_));
 sky130_fd_sc_hd__buf_4 _14947_ (.A(\top_inst.grid_inst.data_path_wires[6][4] ),
    .X(_07615_));
 sky130_fd_sc_hd__nand2_1 _14948_ (.A(_04865_),
    .B(_07378_),
    .Y(_07616_));
 sky130_fd_sc_hd__buf_4 _14949_ (.A(_04868_),
    .X(_07617_));
 sky130_fd_sc_hd__buf_2 _14950_ (.A(_07617_),
    .X(_07618_));
 sky130_fd_sc_hd__o211a_1 _14951_ (.A1(_07615_),
    .A2(_07611_),
    .B1(_07616_),
    .C1(_07618_),
    .X(_00454_));
 sky130_fd_sc_hd__buf_4 _14952_ (.A(\top_inst.grid_inst.data_path_wires[6][5] ),
    .X(_07619_));
 sky130_fd_sc_hd__nand2_1 _14953_ (.A(_04865_),
    .B(_07416_),
    .Y(_07620_));
 sky130_fd_sc_hd__o211a_1 _14954_ (.A1(_07619_),
    .A2(_07611_),
    .B1(_07620_),
    .C1(_07618_),
    .X(_00455_));
 sky130_fd_sc_hd__buf_2 _14955_ (.A(\top_inst.grid_inst.data_path_wires[6][6] ),
    .X(_07621_));
 sky130_fd_sc_hd__buf_4 _14956_ (.A(_07621_),
    .X(_07622_));
 sky130_fd_sc_hd__nand2_1 _14957_ (.A(_04865_),
    .B(_07460_),
    .Y(_07623_));
 sky130_fd_sc_hd__o211a_1 _14958_ (.A1(_07622_),
    .A2(_07611_),
    .B1(_07623_),
    .C1(_07618_),
    .X(_00456_));
 sky130_fd_sc_hd__clkbuf_4 _14959_ (.A(\top_inst.grid_inst.data_path_wires[6][7] ),
    .X(_07624_));
 sky130_fd_sc_hd__or2_1 _14960_ (.A(_05736_),
    .B(_07090_),
    .X(_07625_));
 sky130_fd_sc_hd__o211a_1 _14961_ (.A1(_07624_),
    .A2(_07611_),
    .B1(_07625_),
    .C1(_07618_),
    .X(_00457_));
 sky130_fd_sc_hd__buf_2 _14962_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[0] ),
    .X(_07626_));
 sky130_fd_sc_hd__buf_2 _14963_ (.A(_07626_),
    .X(_07627_));
 sky130_fd_sc_hd__or2_1 _14964_ (.A(_07627_),
    .B(_07075_),
    .X(_07628_));
 sky130_fd_sc_hd__o211a_1 _14965_ (.A1(_07606_),
    .A2(_06647_),
    .B1(_07628_),
    .C1(_07618_),
    .X(_00458_));
 sky130_fd_sc_hd__clkbuf_4 _14966_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[1] ),
    .X(_07629_));
 sky130_fd_sc_hd__or2_1 _14967_ (.A(_07629_),
    .B(_07075_),
    .X(_07630_));
 sky130_fd_sc_hd__o211a_1 _14968_ (.A1(_07608_),
    .A2(_06647_),
    .B1(_07630_),
    .C1(_07618_),
    .X(_00459_));
 sky130_fd_sc_hd__buf_4 _14969_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[2] ),
    .X(_07631_));
 sky130_fd_sc_hd__or2_1 _14970_ (.A(_07631_),
    .B(_07075_),
    .X(_07632_));
 sky130_fd_sc_hd__o211a_1 _14971_ (.A1(_07610_),
    .A2(_06647_),
    .B1(_07632_),
    .C1(_07618_),
    .X(_00460_));
 sky130_fd_sc_hd__clkbuf_4 _14972_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[3] ),
    .X(_07633_));
 sky130_fd_sc_hd__or2_1 _14973_ (.A(_07633_),
    .B(_07075_),
    .X(_07634_));
 sky130_fd_sc_hd__o211a_1 _14974_ (.A1(_07613_),
    .A2(_06647_),
    .B1(_07634_),
    .C1(_07618_),
    .X(_00461_));
 sky130_fd_sc_hd__clkbuf_4 _14975_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[4] ),
    .X(_07635_));
 sky130_fd_sc_hd__or2_1 _14976_ (.A(_07635_),
    .B(_07075_),
    .X(_07636_));
 sky130_fd_sc_hd__o211a_1 _14977_ (.A1(_07615_),
    .A2(_06647_),
    .B1(_07636_),
    .C1(_07618_),
    .X(_00462_));
 sky130_fd_sc_hd__clkbuf_4 _14978_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[5] ),
    .X(_07637_));
 sky130_fd_sc_hd__or2_1 _14979_ (.A(_07637_),
    .B(_07075_),
    .X(_07638_));
 sky130_fd_sc_hd__o211a_1 _14980_ (.A1(_07619_),
    .A2(_06647_),
    .B1(_07638_),
    .C1(_07618_),
    .X(_00463_));
 sky130_fd_sc_hd__clkbuf_4 _14981_ (.A(_05755_),
    .X(_07639_));
 sky130_fd_sc_hd__buf_2 _14982_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[6] ),
    .X(_07640_));
 sky130_fd_sc_hd__buf_2 _14983_ (.A(_05772_),
    .X(_07641_));
 sky130_fd_sc_hd__or2_1 _14984_ (.A(_07640_),
    .B(_07641_),
    .X(_07642_));
 sky130_fd_sc_hd__clkbuf_4 _14985_ (.A(_07617_),
    .X(_07643_));
 sky130_fd_sc_hd__o211a_1 _14986_ (.A1(_07622_),
    .A2(_07639_),
    .B1(_07642_),
    .C1(_07643_),
    .X(_00464_));
 sky130_fd_sc_hd__or2_1 _14987_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[7] ),
    .B(_07641_),
    .X(_07644_));
 sky130_fd_sc_hd__o211a_1 _14988_ (.A1(_07624_),
    .A2(_07639_),
    .B1(_07644_),
    .C1(_07643_),
    .X(_00465_));
 sky130_fd_sc_hd__and3_1 _14989_ (.A(_07606_),
    .B(_07627_),
    .C(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[0] ),
    .X(_07645_));
 sky130_fd_sc_hd__a21oi_1 _14990_ (.A1(_07606_),
    .A2(_07627_),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[0] ),
    .Y(_07646_));
 sky130_fd_sc_hd__o21ai_1 _14991_ (.A1(_07645_),
    .A2(_07646_),
    .B1(_05336_),
    .Y(_07647_));
 sky130_fd_sc_hd__o211a_1 _14992_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[0] ),
    .A2(_06660_),
    .B1(_07647_),
    .C1(_07643_),
    .X(_00466_));
 sky130_fd_sc_hd__a22o_1 _14993_ (.A1(_07606_),
    .A2(_07629_),
    .B1(_07627_),
    .B2(_07608_),
    .X(_07648_));
 sky130_fd_sc_hd__nand4_2 _14994_ (.A(_07608_),
    .B(_07606_),
    .C(_07629_),
    .D(_07627_),
    .Y(_07649_));
 sky130_fd_sc_hd__nand3_2 _14995_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[1] ),
    .B(_07648_),
    .C(_07649_),
    .Y(_07650_));
 sky130_fd_sc_hd__a21o_1 _14996_ (.A1(_07648_),
    .A2(_07649_),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[1] ),
    .X(_07651_));
 sky130_fd_sc_hd__a21o_1 _14997_ (.A1(_07650_),
    .A2(_07651_),
    .B1(_07645_),
    .X(_07652_));
 sky130_fd_sc_hd__nand3_2 _14998_ (.A(_07645_),
    .B(_07650_),
    .C(_07651_),
    .Y(_07653_));
 sky130_fd_sc_hd__a21o_1 _14999_ (.A1(_07652_),
    .A2(_07653_),
    .B1(_06682_),
    .X(_07654_));
 sky130_fd_sc_hd__o211a_1 _15000_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[1] ),
    .A2(_06660_),
    .B1(_07654_),
    .C1(_07643_),
    .X(_00467_));
 sky130_fd_sc_hd__nand2_1 _15001_ (.A(_07606_),
    .B(_07631_),
    .Y(_07655_));
 sky130_fd_sc_hd__a22o_1 _15002_ (.A1(_07608_),
    .A2(_07629_),
    .B1(_07627_),
    .B2(_07610_),
    .X(_07656_));
 sky130_fd_sc_hd__nand4_1 _15003_ (.A(_07610_),
    .B(_07608_),
    .C(_07629_),
    .D(_07627_),
    .Y(_07657_));
 sky130_fd_sc_hd__nand2_1 _15004_ (.A(_07656_),
    .B(_07657_),
    .Y(_07658_));
 sky130_fd_sc_hd__xor2_1 _15005_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[2] ),
    .B(_07658_),
    .X(_07659_));
 sky130_fd_sc_hd__nand2_1 _15006_ (.A(_07649_),
    .B(_07650_),
    .Y(_07660_));
 sky130_fd_sc_hd__xor2_1 _15007_ (.A(_07659_),
    .B(_07660_),
    .X(_07661_));
 sky130_fd_sc_hd__or2_1 _15008_ (.A(_07655_),
    .B(_07661_),
    .X(_07662_));
 sky130_fd_sc_hd__nand2_1 _15009_ (.A(_07655_),
    .B(_07661_),
    .Y(_07663_));
 sky130_fd_sc_hd__and2_1 _15010_ (.A(_07662_),
    .B(_07663_),
    .X(_07664_));
 sky130_fd_sc_hd__xnor2_1 _15011_ (.A(_07653_),
    .B(_07664_),
    .Y(_07665_));
 sky130_fd_sc_hd__or2_1 _15012_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[2] ),
    .B(_06168_),
    .X(_07666_));
 sky130_fd_sc_hd__o211a_1 _15013_ (.A1(_06848_),
    .A2(_07665_),
    .B1(_07666_),
    .C1(_07643_),
    .X(_00468_));
 sky130_fd_sc_hd__or2b_1 _15014_ (.A(_07653_),
    .B_N(_07664_),
    .X(_07667_));
 sky130_fd_sc_hd__or2b_1 _15015_ (.A(_07659_),
    .B_N(_07660_),
    .X(_07668_));
 sky130_fd_sc_hd__a22o_1 _15016_ (.A1(_07606_),
    .A2(_07633_),
    .B1(_07631_),
    .B2(_07608_),
    .X(_07669_));
 sky130_fd_sc_hd__and3_1 _15017_ (.A(\top_inst.grid_inst.data_path_wires[6][1] ),
    .B(\top_inst.grid_inst.data_path_wires[6][0] ),
    .C(_07633_),
    .X(_07670_));
 sky130_fd_sc_hd__nand2_2 _15018_ (.A(_07631_),
    .B(_07670_),
    .Y(_07671_));
 sky130_fd_sc_hd__nand2_1 _15019_ (.A(_07669_),
    .B(_07671_),
    .Y(_07672_));
 sky130_fd_sc_hd__a22o_1 _15020_ (.A1(_07610_),
    .A2(_07629_),
    .B1(_07627_),
    .B2(_07613_),
    .X(_07673_));
 sky130_fd_sc_hd__nand4_1 _15021_ (.A(_07613_),
    .B(_07610_),
    .C(_07629_),
    .D(_07627_),
    .Y(_07674_));
 sky130_fd_sc_hd__and3_1 _15022_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[3] ),
    .B(_07673_),
    .C(_07674_),
    .X(_07675_));
 sky130_fd_sc_hd__a21oi_1 _15023_ (.A1(_07673_),
    .A2(_07674_),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[3] ),
    .Y(_07676_));
 sky130_fd_sc_hd__or2_1 _15024_ (.A(_07675_),
    .B(_07676_),
    .X(_07677_));
 sky130_fd_sc_hd__a21boi_2 _15025_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[2] ),
    .A2(_07656_),
    .B1_N(_07657_),
    .Y(_07678_));
 sky130_fd_sc_hd__xnor2_1 _15026_ (.A(_07677_),
    .B(_07678_),
    .Y(_07679_));
 sky130_fd_sc_hd__xnor2_1 _15027_ (.A(_07672_),
    .B(_07679_),
    .Y(_07680_));
 sky130_fd_sc_hd__a21o_1 _15028_ (.A1(_07668_),
    .A2(_07662_),
    .B1(_07680_),
    .X(_07681_));
 sky130_fd_sc_hd__inv_2 _15029_ (.A(_07681_),
    .Y(_07682_));
 sky130_fd_sc_hd__and3_1 _15030_ (.A(_07668_),
    .B(_07662_),
    .C(_07680_),
    .X(_07683_));
 sky130_fd_sc_hd__or3_1 _15031_ (.A(_07667_),
    .B(_07682_),
    .C(_07683_),
    .X(_07684_));
 sky130_fd_sc_hd__o21ai_1 _15032_ (.A1(_07682_),
    .A2(_07683_),
    .B1(_07667_),
    .Y(_07685_));
 sky130_fd_sc_hd__and2_1 _15033_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[3] ),
    .B(_05326_),
    .X(_07686_));
 sky130_fd_sc_hd__a31o_1 _15034_ (.A1(_05887_),
    .A2(_07684_),
    .A3(_07685_),
    .B1(_07686_),
    .X(_07687_));
 sky130_fd_sc_hd__and2_1 _15035_ (.A(_07117_),
    .B(_07687_),
    .X(_07688_));
 sky130_fd_sc_hd__clkbuf_1 _15036_ (.A(_07688_),
    .X(_00469_));
 sky130_fd_sc_hd__a22o_1 _15037_ (.A1(\top_inst.grid_inst.data_path_wires[6][3] ),
    .A2(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[1] ),
    .B1(_07626_),
    .B2(\top_inst.grid_inst.data_path_wires[6][4] ),
    .X(_07689_));
 sky130_fd_sc_hd__nand4_1 _15038_ (.A(\top_inst.grid_inst.data_path_wires[6][4] ),
    .B(\top_inst.grid_inst.data_path_wires[6][3] ),
    .C(_07629_),
    .D(_07626_),
    .Y(_07690_));
 sky130_fd_sc_hd__nand2_1 _15039_ (.A(_07689_),
    .B(_07690_),
    .Y(_07691_));
 sky130_fd_sc_hd__xor2_2 _15040_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[4] ),
    .B(_07691_),
    .X(_07692_));
 sky130_fd_sc_hd__xor2_2 _15041_ (.A(_07671_),
    .B(_07692_),
    .X(_07693_));
 sky130_fd_sc_hd__a21bo_1 _15042_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[3] ),
    .A2(_07673_),
    .B1_N(_07674_),
    .X(_07694_));
 sky130_fd_sc_hd__xnor2_2 _15043_ (.A(_07693_),
    .B(_07694_),
    .Y(_07695_));
 sky130_fd_sc_hd__nand2_1 _15044_ (.A(_07610_),
    .B(_07631_),
    .Y(_07696_));
 sky130_fd_sc_hd__a22o_1 _15045_ (.A1(\top_inst.grid_inst.data_path_wires[6][0] ),
    .A2(_07635_),
    .B1(_07633_),
    .B2(\top_inst.grid_inst.data_path_wires[6][1] ),
    .X(_07697_));
 sky130_fd_sc_hd__a21bo_1 _15046_ (.A1(_07635_),
    .A2(_07670_),
    .B1_N(_07697_),
    .X(_07698_));
 sky130_fd_sc_hd__xor2_2 _15047_ (.A(_07696_),
    .B(_07698_),
    .X(_07699_));
 sky130_fd_sc_hd__xor2_2 _15048_ (.A(_07695_),
    .B(_07699_),
    .X(_07700_));
 sky130_fd_sc_hd__or2_1 _15049_ (.A(_07672_),
    .B(_07679_),
    .X(_07701_));
 sky130_fd_sc_hd__o21ai_2 _15050_ (.A1(_07677_),
    .A2(_07678_),
    .B1(_07701_),
    .Y(_07702_));
 sky130_fd_sc_hd__xor2_2 _15051_ (.A(_07700_),
    .B(_07702_),
    .X(_07703_));
 sky130_fd_sc_hd__nand2_1 _15052_ (.A(_07681_),
    .B(_07684_),
    .Y(_07704_));
 sky130_fd_sc_hd__nor2_1 _15053_ (.A(_07703_),
    .B(_07704_),
    .Y(_07705_));
 sky130_fd_sc_hd__a21o_1 _15054_ (.A1(_07703_),
    .A2(_07704_),
    .B1(_07057_),
    .X(_07706_));
 sky130_fd_sc_hd__buf_4 _15055_ (.A(_04873_),
    .X(_07707_));
 sky130_fd_sc_hd__clkbuf_8 _15056_ (.A(_07707_),
    .X(_07708_));
 sky130_fd_sc_hd__o221a_1 _15057_ (.A1(net1071),
    .A2(_07048_),
    .B1(_07705_),
    .B2(_07706_),
    .C1(_07708_),
    .X(_00470_));
 sky130_fd_sc_hd__nor2_1 _15058_ (.A(_07684_),
    .B(_07703_),
    .Y(_07709_));
 sky130_fd_sc_hd__and2b_1 _15059_ (.A_N(_07695_),
    .B(_07699_),
    .X(_07710_));
 sky130_fd_sc_hd__nand2_1 _15060_ (.A(_07606_),
    .B(_07637_),
    .Y(_07711_));
 sky130_fd_sc_hd__a22o_1 _15061_ (.A1(\top_inst.grid_inst.data_path_wires[6][1] ),
    .A2(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[6][2] ),
    .X(_07712_));
 sky130_fd_sc_hd__nand4_4 _15062_ (.A(\top_inst.grid_inst.data_path_wires[6][2] ),
    .B(\top_inst.grid_inst.data_path_wires[6][1] ),
    .C(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[3] ),
    .Y(_07713_));
 sky130_fd_sc_hd__a22o_1 _15063_ (.A1(_07613_),
    .A2(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[2] ),
    .B1(_07712_),
    .B2(_07713_),
    .X(_07714_));
 sky130_fd_sc_hd__nand4_2 _15064_ (.A(_07613_),
    .B(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[2] ),
    .C(_07712_),
    .D(_07713_),
    .Y(_07715_));
 sky130_fd_sc_hd__nand2_1 _15065_ (.A(_07714_),
    .B(_07715_),
    .Y(_07716_));
 sky130_fd_sc_hd__or2_1 _15066_ (.A(_07711_),
    .B(_07716_),
    .X(_07717_));
 sky130_fd_sc_hd__nand2_1 _15067_ (.A(_07711_),
    .B(_07716_),
    .Y(_07718_));
 sky130_fd_sc_hd__and2_1 _15068_ (.A(_07717_),
    .B(_07718_),
    .X(_07719_));
 sky130_fd_sc_hd__a21boi_2 _15069_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[4] ),
    .A2(_07689_),
    .B1_N(_07690_),
    .Y(_07720_));
 sky130_fd_sc_hd__a32o_1 _15070_ (.A1(_07610_),
    .A2(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[2] ),
    .A3(_07697_),
    .B1(_07670_),
    .B2(_07635_),
    .X(_07721_));
 sky130_fd_sc_hd__a22o_1 _15071_ (.A1(\top_inst.grid_inst.data_path_wires[6][4] ),
    .A2(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[1] ),
    .B1(_07626_),
    .B2(\top_inst.grid_inst.data_path_wires[6][5] ),
    .X(_07722_));
 sky130_fd_sc_hd__nand4_1 _15072_ (.A(\top_inst.grid_inst.data_path_wires[6][5] ),
    .B(\top_inst.grid_inst.data_path_wires[6][4] ),
    .C(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[1] ),
    .D(_07626_),
    .Y(_07723_));
 sky130_fd_sc_hd__nand2_1 _15073_ (.A(_07722_),
    .B(_07723_),
    .Y(_07724_));
 sky130_fd_sc_hd__xor2_2 _15074_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[5] ),
    .B(_07724_),
    .X(_07725_));
 sky130_fd_sc_hd__xnor2_2 _15075_ (.A(_07721_),
    .B(_07725_),
    .Y(_07726_));
 sky130_fd_sc_hd__xnor2_2 _15076_ (.A(_07720_),
    .B(_07726_),
    .Y(_07727_));
 sky130_fd_sc_hd__xor2_2 _15077_ (.A(_07719_),
    .B(_07727_),
    .X(_07728_));
 sky130_fd_sc_hd__xor2_2 _15078_ (.A(_07710_),
    .B(_07728_),
    .X(_07729_));
 sky130_fd_sc_hd__nor2_1 _15079_ (.A(_07671_),
    .B(_07692_),
    .Y(_07730_));
 sky130_fd_sc_hd__a21o_1 _15080_ (.A1(_07693_),
    .A2(_07694_),
    .B1(_07730_),
    .X(_07731_));
 sky130_fd_sc_hd__xnor2_2 _15081_ (.A(_07729_),
    .B(_07731_),
    .Y(_07732_));
 sky130_fd_sc_hd__or2b_1 _15082_ (.A(_07700_),
    .B_N(_07702_),
    .X(_07733_));
 sky130_fd_sc_hd__o21a_1 _15083_ (.A1(_07681_),
    .A2(_07703_),
    .B1(_07733_),
    .X(_07734_));
 sky130_fd_sc_hd__xor2_1 _15084_ (.A(_07732_),
    .B(_07734_),
    .X(_07735_));
 sky130_fd_sc_hd__nand2_1 _15085_ (.A(_07709_),
    .B(_07735_),
    .Y(_07736_));
 sky130_fd_sc_hd__o21a_1 _15086_ (.A1(_07709_),
    .A2(_07735_),
    .B1(_05315_),
    .X(_07737_));
 sky130_fd_sc_hd__a22o_1 _15087_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[5] ),
    .A2(_06242_),
    .B1(_07736_),
    .B2(_07737_),
    .X(_07738_));
 sky130_fd_sc_hd__and2_1 _15088_ (.A(_07117_),
    .B(_07738_),
    .X(_07739_));
 sky130_fd_sc_hd__clkbuf_1 _15089_ (.A(_07739_),
    .X(_00471_));
 sky130_fd_sc_hd__nor2_1 _15090_ (.A(_07733_),
    .B(_07732_),
    .Y(_07740_));
 sky130_fd_sc_hd__nand2_1 _15091_ (.A(_07710_),
    .B(_07728_),
    .Y(_07741_));
 sky130_fd_sc_hd__nand2_1 _15092_ (.A(_07729_),
    .B(_07731_),
    .Y(_07742_));
 sky130_fd_sc_hd__or2b_1 _15093_ (.A(_07725_),
    .B_N(_07721_),
    .X(_07743_));
 sky130_fd_sc_hd__or2b_1 _15094_ (.A(_07720_),
    .B_N(_07726_),
    .X(_07744_));
 sky130_fd_sc_hd__a22o_1 _15095_ (.A1(\top_inst.grid_inst.data_path_wires[6][0] ),
    .A2(_07640_),
    .B1(_07637_),
    .B2(_07608_),
    .X(_07745_));
 sky130_fd_sc_hd__nand4_2 _15096_ (.A(_07608_),
    .B(\top_inst.grid_inst.data_path_wires[6][0] ),
    .C(_07640_),
    .D(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[5] ),
    .Y(_07746_));
 sky130_fd_sc_hd__nand2_1 _15097_ (.A(_07745_),
    .B(_07746_),
    .Y(_07747_));
 sky130_fd_sc_hd__a22o_1 _15098_ (.A1(\top_inst.grid_inst.data_path_wires[6][2] ),
    .A2(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[6][3] ),
    .X(_07748_));
 sky130_fd_sc_hd__nand4_4 _15099_ (.A(\top_inst.grid_inst.data_path_wires[6][3] ),
    .B(_07610_),
    .C(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[3] ),
    .Y(_07749_));
 sky130_fd_sc_hd__a22o_1 _15100_ (.A1(_07615_),
    .A2(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[2] ),
    .B1(_07748_),
    .B2(_07749_),
    .X(_07750_));
 sky130_fd_sc_hd__nand4_2 _15101_ (.A(_07615_),
    .B(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[2] ),
    .C(_07748_),
    .D(_07749_),
    .Y(_07751_));
 sky130_fd_sc_hd__nand2_1 _15102_ (.A(_07750_),
    .B(_07751_),
    .Y(_07752_));
 sky130_fd_sc_hd__xnor2_1 _15103_ (.A(_07747_),
    .B(_07752_),
    .Y(_07753_));
 sky130_fd_sc_hd__xor2_1 _15104_ (.A(_07717_),
    .B(_07753_),
    .X(_07754_));
 sky130_fd_sc_hd__a21boi_2 _15105_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[5] ),
    .A2(_07722_),
    .B1_N(_07723_),
    .Y(_07755_));
 sky130_fd_sc_hd__a22o_1 _15106_ (.A1(\top_inst.grid_inst.data_path_wires[6][5] ),
    .A2(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[1] ),
    .B1(_07626_),
    .B2(\top_inst.grid_inst.data_path_wires[6][6] ),
    .X(_07756_));
 sky130_fd_sc_hd__nand4_1 _15107_ (.A(_07621_),
    .B(\top_inst.grid_inst.data_path_wires[6][5] ),
    .C(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[1] ),
    .D(_07626_),
    .Y(_07757_));
 sky130_fd_sc_hd__and3_1 _15108_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[6] ),
    .B(_07756_),
    .C(_07757_),
    .X(_07758_));
 sky130_fd_sc_hd__a21oi_1 _15109_ (.A1(_07756_),
    .A2(_07757_),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[6] ),
    .Y(_07759_));
 sky130_fd_sc_hd__a211o_1 _15110_ (.A1(_07713_),
    .A2(_07715_),
    .B1(_07758_),
    .C1(_07759_),
    .X(_07760_));
 sky130_fd_sc_hd__o211ai_1 _15111_ (.A1(_07758_),
    .A2(_07759_),
    .B1(_07713_),
    .C1(_07715_),
    .Y(_07761_));
 sky130_fd_sc_hd__and2_1 _15112_ (.A(_07760_),
    .B(_07761_),
    .X(_07762_));
 sky130_fd_sc_hd__xnor2_1 _15113_ (.A(_07755_),
    .B(_07762_),
    .Y(_07763_));
 sky130_fd_sc_hd__nand2_1 _15114_ (.A(_07754_),
    .B(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__or2_1 _15115_ (.A(_07754_),
    .B(_07763_),
    .X(_07765_));
 sky130_fd_sc_hd__and2_1 _15116_ (.A(_07719_),
    .B(_07727_),
    .X(_07766_));
 sky130_fd_sc_hd__a21oi_1 _15117_ (.A1(_07764_),
    .A2(_07765_),
    .B1(_07766_),
    .Y(_07767_));
 sky130_fd_sc_hd__and3_1 _15118_ (.A(_07766_),
    .B(_07764_),
    .C(_07765_),
    .X(_07768_));
 sky130_fd_sc_hd__a211oi_2 _15119_ (.A1(_07743_),
    .A2(_07744_),
    .B1(_07767_),
    .C1(_07768_),
    .Y(_07769_));
 sky130_fd_sc_hd__o211a_1 _15120_ (.A1(_07767_),
    .A2(_07768_),
    .B1(_07743_),
    .C1(_07744_),
    .X(_07770_));
 sky130_fd_sc_hd__a211o_1 _15121_ (.A1(_07741_),
    .A2(_07742_),
    .B1(_07769_),
    .C1(_07770_),
    .X(_07771_));
 sky130_fd_sc_hd__o211ai_1 _15122_ (.A1(_07769_),
    .A2(_07770_),
    .B1(_07741_),
    .C1(_07742_),
    .Y(_07772_));
 sky130_fd_sc_hd__and3_1 _15123_ (.A(_07740_),
    .B(_07771_),
    .C(_07772_),
    .X(_07773_));
 sky130_fd_sc_hd__a21oi_1 _15124_ (.A1(_07771_),
    .A2(_07772_),
    .B1(_07740_),
    .Y(_07774_));
 sky130_fd_sc_hd__nor2_1 _15125_ (.A(_07773_),
    .B(_07774_),
    .Y(_07775_));
 sky130_fd_sc_hd__o31a_1 _15126_ (.A1(_07681_),
    .A2(_07703_),
    .A3(_07732_),
    .B1(_07736_),
    .X(_07776_));
 sky130_fd_sc_hd__xnor2_1 _15127_ (.A(_07775_),
    .B(_07776_),
    .Y(_07777_));
 sky130_fd_sc_hd__mux2_1 _15128_ (.A0(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[6] ),
    .A1(_07777_),
    .S(_06701_),
    .X(_07778_));
 sky130_fd_sc_hd__and2_1 _15129_ (.A(_07117_),
    .B(_07778_),
    .X(_07779_));
 sky130_fd_sc_hd__clkbuf_1 _15130_ (.A(_07779_),
    .X(_00472_));
 sky130_fd_sc_hd__nor2_1 _15131_ (.A(_07747_),
    .B(_07752_),
    .Y(_07780_));
 sky130_fd_sc_hd__nand2_1 _15132_ (.A(\top_inst.grid_inst.data_path_wires[6][1] ),
    .B(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[6] ),
    .Y(_07781_));
 sky130_fd_sc_hd__or2b_1 _15133_ (.A(\top_inst.grid_inst.data_path_wires[6][0] ),
    .B_N(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[7] ),
    .X(_07782_));
 sky130_fd_sc_hd__xnor2_1 _15134_ (.A(_07781_),
    .B(_07782_),
    .Y(_07783_));
 sky130_fd_sc_hd__nand2_1 _15135_ (.A(\top_inst.grid_inst.data_path_wires[6][2] ),
    .B(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[5] ),
    .Y(_07784_));
 sky130_fd_sc_hd__xnor2_1 _15136_ (.A(_07783_),
    .B(_07784_),
    .Y(_07785_));
 sky130_fd_sc_hd__xor2_1 _15137_ (.A(_07746_),
    .B(_07785_),
    .X(_07786_));
 sky130_fd_sc_hd__a22o_1 _15138_ (.A1(\top_inst.grid_inst.data_path_wires[6][3] ),
    .A2(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[6][4] ),
    .X(_07787_));
 sky130_fd_sc_hd__nand4_2 _15139_ (.A(\top_inst.grid_inst.data_path_wires[6][4] ),
    .B(\top_inst.grid_inst.data_path_wires[6][3] ),
    .C(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[3] ),
    .Y(_07788_));
 sky130_fd_sc_hd__a22o_1 _15140_ (.A1(_07619_),
    .A2(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[2] ),
    .B1(_07787_),
    .B2(_07788_),
    .X(_07789_));
 sky130_fd_sc_hd__nand4_2 _15141_ (.A(_07619_),
    .B(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[2] ),
    .C(_07787_),
    .D(_07788_),
    .Y(_07790_));
 sky130_fd_sc_hd__nand2_1 _15142_ (.A(_07789_),
    .B(_07790_),
    .Y(_07791_));
 sky130_fd_sc_hd__xnor2_1 _15143_ (.A(_07786_),
    .B(_07791_),
    .Y(_07792_));
 sky130_fd_sc_hd__xnor2_1 _15144_ (.A(_07780_),
    .B(_07792_),
    .Y(_07793_));
 sky130_fd_sc_hd__a21bo_1 _15145_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[6] ),
    .A2(_07756_),
    .B1_N(_07757_),
    .X(_07794_));
 sky130_fd_sc_hd__a22o_1 _15146_ (.A1(_07621_),
    .A2(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[1] ),
    .B1(_07626_),
    .B2(\top_inst.grid_inst.data_path_wires[6][7] ),
    .X(_07795_));
 sky130_fd_sc_hd__nand4_1 _15147_ (.A(\top_inst.grid_inst.data_path_wires[6][7] ),
    .B(_07621_),
    .C(_07629_),
    .D(_07626_),
    .Y(_07796_));
 sky130_fd_sc_hd__and3_1 _15148_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[7] ),
    .B(_07795_),
    .C(_07796_),
    .X(_07797_));
 sky130_fd_sc_hd__a21oi_1 _15149_ (.A1(_07795_),
    .A2(_07796_),
    .B1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[7] ),
    .Y(_07798_));
 sky130_fd_sc_hd__a211oi_2 _15150_ (.A1(_07749_),
    .A2(_07751_),
    .B1(_07797_),
    .C1(_07798_),
    .Y(_07799_));
 sky130_fd_sc_hd__o211a_1 _15151_ (.A1(_07797_),
    .A2(_07798_),
    .B1(_07749_),
    .C1(_07751_),
    .X(_07800_));
 sky130_fd_sc_hd__nor2_1 _15152_ (.A(_07799_),
    .B(_07800_),
    .Y(_07801_));
 sky130_fd_sc_hd__xnor2_1 _15153_ (.A(_07794_),
    .B(_07801_),
    .Y(_07802_));
 sky130_fd_sc_hd__xor2_1 _15154_ (.A(_07793_),
    .B(_07802_),
    .X(_07803_));
 sky130_fd_sc_hd__o21ai_1 _15155_ (.A1(_07717_),
    .A2(_07753_),
    .B1(_07764_),
    .Y(_07804_));
 sky130_fd_sc_hd__xnor2_1 _15156_ (.A(_07803_),
    .B(_07804_),
    .Y(_07805_));
 sky130_fd_sc_hd__or2b_1 _15157_ (.A(_07755_),
    .B_N(_07762_),
    .X(_07806_));
 sky130_fd_sc_hd__nand2_1 _15158_ (.A(_07760_),
    .B(_07806_),
    .Y(_07807_));
 sky130_fd_sc_hd__xnor2_1 _15159_ (.A(_07805_),
    .B(_07807_),
    .Y(_07808_));
 sky130_fd_sc_hd__nor2_1 _15160_ (.A(_07768_),
    .B(_07769_),
    .Y(_07809_));
 sky130_fd_sc_hd__xnor2_1 _15161_ (.A(_07808_),
    .B(_07809_),
    .Y(_07810_));
 sky130_fd_sc_hd__xnor2_1 _15162_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[7] ),
    .B(_07810_),
    .Y(_07811_));
 sky130_fd_sc_hd__xor2_1 _15163_ (.A(_07771_),
    .B(_07811_),
    .X(_07812_));
 sky130_fd_sc_hd__o21bai_1 _15164_ (.A1(_07774_),
    .A2(_07776_),
    .B1_N(_07773_),
    .Y(_07813_));
 sky130_fd_sc_hd__nor2_1 _15165_ (.A(_07812_),
    .B(_07813_),
    .Y(_07814_));
 sky130_fd_sc_hd__a21o_1 _15166_ (.A1(_07812_),
    .A2(_07813_),
    .B1(_06404_),
    .X(_07815_));
 sky130_fd_sc_hd__buf_6 _15167_ (.A(_05326_),
    .X(_07816_));
 sky130_fd_sc_hd__a2bb2o_1 _15168_ (.A1_N(_07814_),
    .A2_N(_07815_),
    .B1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[7] ),
    .B2(_07816_),
    .X(_07817_));
 sky130_fd_sc_hd__and2_1 _15169_ (.A(_07117_),
    .B(_07817_),
    .X(_07818_));
 sky130_fd_sc_hd__clkbuf_1 _15170_ (.A(_07818_),
    .X(_00473_));
 sky130_fd_sc_hd__nor2_1 _15171_ (.A(_07771_),
    .B(_07811_),
    .Y(_07819_));
 sky130_fd_sc_hd__a21o_1 _15172_ (.A1(_07812_),
    .A2(_07813_),
    .B1(_07819_),
    .X(_07820_));
 sky130_fd_sc_hd__or2b_1 _15173_ (.A(_07809_),
    .B_N(_07808_),
    .X(_07821_));
 sky130_fd_sc_hd__nand2_1 _15174_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[7] ),
    .B(_07810_),
    .Y(_07822_));
 sky130_fd_sc_hd__and4b_1 _15175_ (.A_N(\top_inst.grid_inst.data_path_wires[6][1] ),
    .B(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[7] ),
    .C(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[6] ),
    .D(\top_inst.grid_inst.data_path_wires[6][2] ),
    .X(_07823_));
 sky130_fd_sc_hd__inv_2 _15176_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[7] ),
    .Y(_07824_));
 sky130_fd_sc_hd__o2bb2a_1 _15177_ (.A1_N(\top_inst.grid_inst.data_path_wires[6][2] ),
    .A2_N(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[6] ),
    .B1(_07824_),
    .B2(\top_inst.grid_inst.data_path_wires[6][1] ),
    .X(_07825_));
 sky130_fd_sc_hd__nor2_1 _15178_ (.A(_07823_),
    .B(_07825_),
    .Y(_07826_));
 sky130_fd_sc_hd__nand2_1 _15179_ (.A(_07613_),
    .B(_07637_),
    .Y(_07827_));
 sky130_fd_sc_hd__xnor2_2 _15180_ (.A(_07826_),
    .B(_07827_),
    .Y(_07828_));
 sky130_fd_sc_hd__nor2_1 _15181_ (.A(_07783_),
    .B(_07784_),
    .Y(_07829_));
 sky130_fd_sc_hd__o21ba_1 _15182_ (.A1(_07781_),
    .A2(_07782_),
    .B1_N(_07829_),
    .X(_07830_));
 sky130_fd_sc_hd__xnor2_2 _15183_ (.A(_07828_),
    .B(_07830_),
    .Y(_07831_));
 sky130_fd_sc_hd__a22o_1 _15184_ (.A1(_07615_),
    .A2(_07635_),
    .B1(_07633_),
    .B2(_07619_),
    .X(_07832_));
 sky130_fd_sc_hd__nand4_4 _15185_ (.A(_07619_),
    .B(_07615_),
    .C(_07635_),
    .D(_07633_),
    .Y(_07833_));
 sky130_fd_sc_hd__a22o_1 _15186_ (.A1(_07621_),
    .A2(_07631_),
    .B1(_07832_),
    .B2(_07833_),
    .X(_07834_));
 sky130_fd_sc_hd__nand4_4 _15187_ (.A(_07622_),
    .B(_07631_),
    .C(_07832_),
    .D(_07833_),
    .Y(_07835_));
 sky130_fd_sc_hd__nand2_1 _15188_ (.A(_07834_),
    .B(_07835_),
    .Y(_07836_));
 sky130_fd_sc_hd__xnor2_1 _15189_ (.A(_07831_),
    .B(_07836_),
    .Y(_07837_));
 sky130_fd_sc_hd__and3_1 _15190_ (.A(_07786_),
    .B(_07789_),
    .C(_07790_),
    .X(_07838_));
 sky130_fd_sc_hd__o21ba_1 _15191_ (.A1(_07746_),
    .A2(_07785_),
    .B1_N(_07838_),
    .X(_07839_));
 sky130_fd_sc_hd__xnor2_1 _15192_ (.A(_07837_),
    .B(_07839_),
    .Y(_07840_));
 sky130_fd_sc_hd__and4_1 _15193_ (.A(_07624_),
    .B(_07622_),
    .C(_07629_),
    .D(_07627_),
    .X(_07841_));
 sky130_fd_sc_hd__o21ai_1 _15194_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[1] ),
    .A2(_07626_),
    .B1(\top_inst.grid_inst.data_path_wires[6][7] ),
    .Y(_07842_));
 sky130_fd_sc_hd__and3_1 _15195_ (.A(\top_inst.grid_inst.data_path_wires[6][7] ),
    .B(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[1] ),
    .C(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[0] ),
    .X(_07843_));
 sky130_fd_sc_hd__clkbuf_4 _15196_ (.A(_07843_),
    .X(_07844_));
 sky130_fd_sc_hd__nor2_4 _15197_ (.A(_07842_),
    .B(_07844_),
    .Y(_07845_));
 sky130_fd_sc_hd__xnor2_1 _15198_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[8] ),
    .B(_07845_),
    .Y(_07846_));
 sky130_fd_sc_hd__a21oi_1 _15199_ (.A1(_07788_),
    .A2(_07790_),
    .B1(_07846_),
    .Y(_07847_));
 sky130_fd_sc_hd__and3_1 _15200_ (.A(_07788_),
    .B(_07790_),
    .C(_07846_),
    .X(_07848_));
 sky130_fd_sc_hd__nor2_1 _15201_ (.A(_07847_),
    .B(_07848_),
    .Y(_07849_));
 sky130_fd_sc_hd__o21a_1 _15202_ (.A1(_07841_),
    .A2(_07797_),
    .B1(_07849_),
    .X(_07850_));
 sky130_fd_sc_hd__nor3_1 _15203_ (.A(_07841_),
    .B(_07797_),
    .C(_07849_),
    .Y(_07851_));
 sky130_fd_sc_hd__nor2_1 _15204_ (.A(_07850_),
    .B(_07851_),
    .Y(_07852_));
 sky130_fd_sc_hd__xnor2_1 _15205_ (.A(_07840_),
    .B(_07852_),
    .Y(_07853_));
 sky130_fd_sc_hd__nand2_1 _15206_ (.A(_07780_),
    .B(_07792_),
    .Y(_07854_));
 sky130_fd_sc_hd__o21a_1 _15207_ (.A1(_07793_),
    .A2(_07802_),
    .B1(_07854_),
    .X(_07855_));
 sky130_fd_sc_hd__xnor2_1 _15208_ (.A(_07853_),
    .B(_07855_),
    .Y(_07856_));
 sky130_fd_sc_hd__a21oi_2 _15209_ (.A1(_07794_),
    .A2(_07801_),
    .B1(_07799_),
    .Y(_07857_));
 sky130_fd_sc_hd__xnor2_1 _15210_ (.A(_07856_),
    .B(_07857_),
    .Y(_07858_));
 sky130_fd_sc_hd__and2b_1 _15211_ (.A_N(_07805_),
    .B(_07807_),
    .X(_07859_));
 sky130_fd_sc_hd__a21oi_1 _15212_ (.A1(_07803_),
    .A2(_07804_),
    .B1(_07859_),
    .Y(_07860_));
 sky130_fd_sc_hd__xnor2_1 _15213_ (.A(_07858_),
    .B(_07860_),
    .Y(_07861_));
 sky130_fd_sc_hd__a21o_1 _15214_ (.A1(_07821_),
    .A2(_07822_),
    .B1(_07861_),
    .X(_07862_));
 sky130_fd_sc_hd__nand3_1 _15215_ (.A(_07821_),
    .B(_07822_),
    .C(_07861_),
    .Y(_07863_));
 sky130_fd_sc_hd__and2_1 _15216_ (.A(_07862_),
    .B(_07863_),
    .X(_07864_));
 sky130_fd_sc_hd__xor2_1 _15217_ (.A(_07820_),
    .B(_07864_),
    .X(_07865_));
 sky130_fd_sc_hd__clkbuf_4 _15218_ (.A(_05312_),
    .X(_07866_));
 sky130_fd_sc_hd__or2_1 _15219_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[8] ),
    .B(_07866_),
    .X(_07867_));
 sky130_fd_sc_hd__o211a_1 _15220_ (.A1(_06848_),
    .A2(_07865_),
    .B1(_07867_),
    .C1(_07643_),
    .X(_00474_));
 sky130_fd_sc_hd__a21bo_1 _15221_ (.A1(_07820_),
    .A2(_07864_),
    .B1_N(_07862_),
    .X(_07868_));
 sky130_fd_sc_hd__or2_1 _15222_ (.A(_07858_),
    .B(_07860_),
    .X(_07869_));
 sky130_fd_sc_hd__and4b_1 _15223_ (.A_N(\top_inst.grid_inst.data_path_wires[6][2] ),
    .B(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[7] ),
    .C(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[6] ),
    .D(\top_inst.grid_inst.data_path_wires[6][3] ),
    .X(_07870_));
 sky130_fd_sc_hd__o2bb2a_1 _15224_ (.A1_N(\top_inst.grid_inst.data_path_wires[6][3] ),
    .A2_N(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[6] ),
    .B1(_07824_),
    .B2(\top_inst.grid_inst.data_path_wires[6][2] ),
    .X(_07871_));
 sky130_fd_sc_hd__nor2_1 _15225_ (.A(_07870_),
    .B(_07871_),
    .Y(_07872_));
 sky130_fd_sc_hd__nand2_1 _15226_ (.A(_07615_),
    .B(_07637_),
    .Y(_07873_));
 sky130_fd_sc_hd__xnor2_1 _15227_ (.A(_07872_),
    .B(_07873_),
    .Y(_07874_));
 sky130_fd_sc_hd__o21ba_1 _15228_ (.A1(_07825_),
    .A2(_07827_),
    .B1_N(_07823_),
    .X(_07875_));
 sky130_fd_sc_hd__xor2_1 _15229_ (.A(_07874_),
    .B(_07875_),
    .X(_07876_));
 sky130_fd_sc_hd__a22o_1 _15230_ (.A1(_07619_),
    .A2(_07635_),
    .B1(_07633_),
    .B2(_07621_),
    .X(_07877_));
 sky130_fd_sc_hd__and4_1 _15231_ (.A(\top_inst.grid_inst.data_path_wires[6][6] ),
    .B(\top_inst.grid_inst.data_path_wires[6][5] ),
    .C(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[3] ),
    .X(_07878_));
 sky130_fd_sc_hd__inv_2 _15232_ (.A(_07878_),
    .Y(_07879_));
 sky130_fd_sc_hd__and2_1 _15233_ (.A(_07877_),
    .B(_07879_),
    .X(_07880_));
 sky130_fd_sc_hd__nand2_4 _15234_ (.A(\top_inst.grid_inst.data_path_wires[6][7] ),
    .B(_07631_),
    .Y(_07881_));
 sky130_fd_sc_hd__xor2_1 _15235_ (.A(_07880_),
    .B(_07881_),
    .X(_07882_));
 sky130_fd_sc_hd__xor2_1 _15236_ (.A(_07876_),
    .B(_07882_),
    .X(_07883_));
 sky130_fd_sc_hd__inv_2 _15237_ (.A(_07830_),
    .Y(_07884_));
 sky130_fd_sc_hd__a32oi_4 _15238_ (.A1(_07831_),
    .A2(_07834_),
    .A3(_07835_),
    .B1(_07884_),
    .B2(_07828_),
    .Y(_07885_));
 sky130_fd_sc_hd__xnor2_1 _15239_ (.A(_07883_),
    .B(_07885_),
    .Y(_07886_));
 sky130_fd_sc_hd__a21o_1 _15240_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[8] ),
    .A2(_07845_),
    .B1(_07844_),
    .X(_07887_));
 sky130_fd_sc_hd__xnor2_1 _15241_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[9] ),
    .B(_07845_),
    .Y(_07888_));
 sky130_fd_sc_hd__a21oi_1 _15242_ (.A1(_07833_),
    .A2(_07835_),
    .B1(_07888_),
    .Y(_07889_));
 sky130_fd_sc_hd__and3_1 _15243_ (.A(_07833_),
    .B(_07835_),
    .C(_07888_),
    .X(_07890_));
 sky130_fd_sc_hd__nor2_1 _15244_ (.A(_07889_),
    .B(_07890_),
    .Y(_07891_));
 sky130_fd_sc_hd__xor2_2 _15245_ (.A(_07887_),
    .B(_07891_),
    .X(_07892_));
 sky130_fd_sc_hd__xnor2_1 _15246_ (.A(_07886_),
    .B(_07892_),
    .Y(_07893_));
 sky130_fd_sc_hd__and2b_1 _15247_ (.A_N(_07839_),
    .B(_07837_),
    .X(_07894_));
 sky130_fd_sc_hd__a21oi_1 _15248_ (.A1(_07840_),
    .A2(_07852_),
    .B1(_07894_),
    .Y(_07895_));
 sky130_fd_sc_hd__xnor2_1 _15249_ (.A(_07893_),
    .B(_07895_),
    .Y(_07896_));
 sky130_fd_sc_hd__nor2_1 _15250_ (.A(_07847_),
    .B(_07850_),
    .Y(_07897_));
 sky130_fd_sc_hd__xnor2_1 _15251_ (.A(_07896_),
    .B(_07897_),
    .Y(_07898_));
 sky130_fd_sc_hd__or2_1 _15252_ (.A(_07853_),
    .B(_07855_),
    .X(_07899_));
 sky130_fd_sc_hd__o21a_1 _15253_ (.A1(_07856_),
    .A2(_07857_),
    .B1(_07899_),
    .X(_07900_));
 sky130_fd_sc_hd__nor2_1 _15254_ (.A(_07898_),
    .B(_07900_),
    .Y(_07901_));
 sky130_fd_sc_hd__and2_1 _15255_ (.A(_07898_),
    .B(_07900_),
    .X(_07902_));
 sky130_fd_sc_hd__or2_1 _15256_ (.A(_07901_),
    .B(_07902_),
    .X(_07903_));
 sky130_fd_sc_hd__xor2_1 _15257_ (.A(_07869_),
    .B(_07903_),
    .X(_07904_));
 sky130_fd_sc_hd__xor2_1 _15258_ (.A(_07868_),
    .B(_07904_),
    .X(_07905_));
 sky130_fd_sc_hd__or2_1 _15259_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[9] ),
    .B(_07866_),
    .X(_07906_));
 sky130_fd_sc_hd__o211a_1 _15260_ (.A1(_06848_),
    .A2(_07905_),
    .B1(_07906_),
    .C1(_07643_),
    .X(_00475_));
 sky130_fd_sc_hd__or2b_1 _15261_ (.A(_07875_),
    .B_N(_07874_),
    .X(_07907_));
 sky130_fd_sc_hd__o21a_1 _15262_ (.A1(_07876_),
    .A2(_07882_),
    .B1(_07907_),
    .X(_07908_));
 sky130_fd_sc_hd__and4b_1 _15263_ (.A_N(_07613_),
    .B(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[7] ),
    .C(_07640_),
    .D(_07615_),
    .X(_07909_));
 sky130_fd_sc_hd__o2bb2a_1 _15264_ (.A1_N(_07615_),
    .A2_N(_07640_),
    .B1(_07824_),
    .B2(_07613_),
    .X(_07910_));
 sky130_fd_sc_hd__nor2_1 _15265_ (.A(_07909_),
    .B(_07910_),
    .Y(_07911_));
 sky130_fd_sc_hd__nand2_1 _15266_ (.A(_07619_),
    .B(_07637_),
    .Y(_07912_));
 sky130_fd_sc_hd__xnor2_1 _15267_ (.A(_07911_),
    .B(_07912_),
    .Y(_07913_));
 sky130_fd_sc_hd__o21ba_1 _15268_ (.A1(_07871_),
    .A2(_07873_),
    .B1_N(_07870_),
    .X(_07914_));
 sky130_fd_sc_hd__xnor2_1 _15269_ (.A(_07913_),
    .B(_07914_),
    .Y(_07915_));
 sky130_fd_sc_hd__and3_1 _15270_ (.A(\top_inst.grid_inst.data_path_wires[6][7] ),
    .B(_07635_),
    .C(_07633_),
    .X(_07916_));
 sky130_fd_sc_hd__a22o_1 _15271_ (.A1(_07621_),
    .A2(_07635_),
    .B1(_07633_),
    .B2(\top_inst.grid_inst.data_path_wires[6][7] ),
    .X(_07917_));
 sky130_fd_sc_hd__a21bo_1 _15272_ (.A1(_07622_),
    .A2(_07916_),
    .B1_N(_07917_),
    .X(_07918_));
 sky130_fd_sc_hd__xor2_1 _15273_ (.A(_07881_),
    .B(_07918_),
    .X(_07919_));
 sky130_fd_sc_hd__xor2_1 _15274_ (.A(_07915_),
    .B(_07919_),
    .X(_07920_));
 sky130_fd_sc_hd__and2b_1 _15275_ (.A_N(_07908_),
    .B(_07920_),
    .X(_07921_));
 sky130_fd_sc_hd__and2b_1 _15276_ (.A_N(_07920_),
    .B(_07908_),
    .X(_07922_));
 sky130_fd_sc_hd__nor2_1 _15277_ (.A(_07921_),
    .B(_07922_),
    .Y(_07923_));
 sky130_fd_sc_hd__clkbuf_4 _15278_ (.A(_07845_),
    .X(_07924_));
 sky130_fd_sc_hd__a21o_1 _15279_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[9] ),
    .A2(_07924_),
    .B1(_07844_),
    .X(_07925_));
 sky130_fd_sc_hd__a31o_1 _15280_ (.A1(_07624_),
    .A2(_07631_),
    .A3(_07877_),
    .B1(_07878_),
    .X(_07926_));
 sky130_fd_sc_hd__xnor2_2 _15281_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[10] ),
    .B(_07845_),
    .Y(_07927_));
 sky130_fd_sc_hd__xnor2_2 _15282_ (.A(_07926_),
    .B(_07927_),
    .Y(_07928_));
 sky130_fd_sc_hd__xor2_2 _15283_ (.A(_07925_),
    .B(_07928_),
    .X(_07929_));
 sky130_fd_sc_hd__xnor2_2 _15284_ (.A(_07923_),
    .B(_07929_),
    .Y(_07930_));
 sky130_fd_sc_hd__and2b_1 _15285_ (.A_N(_07885_),
    .B(_07883_),
    .X(_07931_));
 sky130_fd_sc_hd__a21oi_2 _15286_ (.A1(_07886_),
    .A2(_07892_),
    .B1(_07931_),
    .Y(_07932_));
 sky130_fd_sc_hd__xnor2_2 _15287_ (.A(_07930_),
    .B(_07932_),
    .Y(_07933_));
 sky130_fd_sc_hd__a21oi_2 _15288_ (.A1(_07887_),
    .A2(_07891_),
    .B1(_07889_),
    .Y(_07934_));
 sky130_fd_sc_hd__xnor2_2 _15289_ (.A(_07933_),
    .B(_07934_),
    .Y(_07935_));
 sky130_fd_sc_hd__or2_1 _15290_ (.A(_07893_),
    .B(_07895_),
    .X(_07936_));
 sky130_fd_sc_hd__o21a_1 _15291_ (.A1(_07896_),
    .A2(_07897_),
    .B1(_07936_),
    .X(_07937_));
 sky130_fd_sc_hd__xor2_1 _15292_ (.A(_07935_),
    .B(_07937_),
    .X(_07938_));
 sky130_fd_sc_hd__and2_1 _15293_ (.A(_07901_),
    .B(_07938_),
    .X(_07939_));
 sky130_fd_sc_hd__nor2_1 _15294_ (.A(_07901_),
    .B(_07938_),
    .Y(_07940_));
 sky130_fd_sc_hd__nor2_1 _15295_ (.A(_07939_),
    .B(_07940_),
    .Y(_07941_));
 sky130_fd_sc_hd__a21oi_1 _15296_ (.A1(_07869_),
    .A2(_07862_),
    .B1(_07903_),
    .Y(_07942_));
 sky130_fd_sc_hd__a31o_1 _15297_ (.A1(_07820_),
    .A2(_07864_),
    .A3(_07904_),
    .B1(_07942_),
    .X(_07943_));
 sky130_fd_sc_hd__nand2_1 _15298_ (.A(_07941_),
    .B(_07943_),
    .Y(_07944_));
 sky130_fd_sc_hd__o21a_1 _15299_ (.A1(_07941_),
    .A2(_07943_),
    .B1(_05315_),
    .X(_07945_));
 sky130_fd_sc_hd__a22o_1 _15300_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[10] ),
    .A2(_06242_),
    .B1(_07944_),
    .B2(_07945_),
    .X(_07946_));
 sky130_fd_sc_hd__and2_1 _15301_ (.A(_07117_),
    .B(_07946_),
    .X(_07947_));
 sky130_fd_sc_hd__clkbuf_1 _15302_ (.A(_07947_),
    .X(_00476_));
 sky130_fd_sc_hd__inv_2 _15303_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[11] ),
    .Y(_07948_));
 sky130_fd_sc_hd__nor2_1 _15304_ (.A(_07935_),
    .B(_07937_),
    .Y(_07949_));
 sky130_fd_sc_hd__nor2_1 _15305_ (.A(_07930_),
    .B(_07932_),
    .Y(_07950_));
 sky130_fd_sc_hd__nor2_1 _15306_ (.A(_07933_),
    .B(_07934_),
    .Y(_07951_));
 sky130_fd_sc_hd__or2b_1 _15307_ (.A(_07914_),
    .B_N(_07913_),
    .X(_07952_));
 sky130_fd_sc_hd__nand2_1 _15308_ (.A(_07915_),
    .B(_07919_),
    .Y(_07953_));
 sky130_fd_sc_hd__o21ai_1 _15309_ (.A1(_07635_),
    .A2(_07633_),
    .B1(\top_inst.grid_inst.data_path_wires[6][7] ),
    .Y(_07954_));
 sky130_fd_sc_hd__nor2_2 _15310_ (.A(_07916_),
    .B(_07954_),
    .Y(_07955_));
 sky130_fd_sc_hd__xnor2_4 _15311_ (.A(_07881_),
    .B(_07955_),
    .Y(_07956_));
 sky130_fd_sc_hd__inv_2 _15312_ (.A(\top_inst.grid_inst.data_path_wires[6][4] ),
    .Y(_07957_));
 sky130_fd_sc_hd__and4_1 _15313_ (.A(\top_inst.grid_inst.data_path_wires[6][5] ),
    .B(_07957_),
    .C(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[7] ),
    .D(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[6] ),
    .X(_07958_));
 sky130_fd_sc_hd__a22o_1 _15314_ (.A1(_07957_),
    .A2(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[7] ),
    .B1(_07640_),
    .B2(\top_inst.grid_inst.data_path_wires[6][5] ),
    .X(_07959_));
 sky130_fd_sc_hd__and2b_1 _15315_ (.A_N(_07958_),
    .B(_07959_),
    .X(_07960_));
 sky130_fd_sc_hd__nand2_1 _15316_ (.A(_07621_),
    .B(_07637_),
    .Y(_07961_));
 sky130_fd_sc_hd__xnor2_1 _15317_ (.A(_07960_),
    .B(_07961_),
    .Y(_07962_));
 sky130_fd_sc_hd__o21ba_1 _15318_ (.A1(_07910_),
    .A2(_07912_),
    .B1_N(_07909_),
    .X(_07963_));
 sky130_fd_sc_hd__xnor2_1 _15319_ (.A(_07962_),
    .B(_07963_),
    .Y(_07964_));
 sky130_fd_sc_hd__nand2_1 _15320_ (.A(_07956_),
    .B(_07964_),
    .Y(_07965_));
 sky130_fd_sc_hd__or2_1 _15321_ (.A(_07956_),
    .B(_07964_),
    .X(_07966_));
 sky130_fd_sc_hd__nand2_1 _15322_ (.A(_07965_),
    .B(_07966_),
    .Y(_07967_));
 sky130_fd_sc_hd__a21oi_1 _15323_ (.A1(_07952_),
    .A2(_07953_),
    .B1(_07967_),
    .Y(_07968_));
 sky130_fd_sc_hd__nand3_1 _15324_ (.A(_07952_),
    .B(_07953_),
    .C(_07967_),
    .Y(_07969_));
 sky130_fd_sc_hd__or2b_1 _15325_ (.A(_07968_),
    .B_N(_07969_),
    .X(_07970_));
 sky130_fd_sc_hd__a21o_1 _15326_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[10] ),
    .A2(_07924_),
    .B1(_07844_),
    .X(_07971_));
 sky130_fd_sc_hd__a32o_1 _15327_ (.A1(_07624_),
    .A2(_07631_),
    .A3(_07917_),
    .B1(_07916_),
    .B2(_07622_),
    .X(_07972_));
 sky130_fd_sc_hd__xnor2_2 _15328_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[11] ),
    .B(_07845_),
    .Y(_07973_));
 sky130_fd_sc_hd__xnor2_2 _15329_ (.A(_07972_),
    .B(_07973_),
    .Y(_07974_));
 sky130_fd_sc_hd__xor2_2 _15330_ (.A(_07971_),
    .B(_07974_),
    .X(_07975_));
 sky130_fd_sc_hd__xnor2_1 _15331_ (.A(_07970_),
    .B(_07975_),
    .Y(_07976_));
 sky130_fd_sc_hd__a21o_1 _15332_ (.A1(_07923_),
    .A2(_07929_),
    .B1(_07921_),
    .X(_07977_));
 sky130_fd_sc_hd__xnor2_1 _15333_ (.A(_07976_),
    .B(_07977_),
    .Y(_07978_));
 sky130_fd_sc_hd__or2b_1 _15334_ (.A(_07927_),
    .B_N(_07926_),
    .X(_07979_));
 sky130_fd_sc_hd__a21bo_1 _15335_ (.A1(_07925_),
    .A2(_07928_),
    .B1_N(_07979_),
    .X(_07980_));
 sky130_fd_sc_hd__xnor2_1 _15336_ (.A(_07978_),
    .B(_07980_),
    .Y(_07981_));
 sky130_fd_sc_hd__o21ai_2 _15337_ (.A1(_07950_),
    .A2(_07951_),
    .B1(_07981_),
    .Y(_07982_));
 sky130_fd_sc_hd__or3_1 _15338_ (.A(_07950_),
    .B(_07951_),
    .C(_07981_),
    .X(_07983_));
 sky130_fd_sc_hd__and2_1 _15339_ (.A(_07982_),
    .B(_07983_),
    .X(_07984_));
 sky130_fd_sc_hd__xnor2_1 _15340_ (.A(_07949_),
    .B(_07984_),
    .Y(_07985_));
 sky130_fd_sc_hd__a21oi_1 _15341_ (.A1(_07941_),
    .A2(_07943_),
    .B1(_07939_),
    .Y(_07986_));
 sky130_fd_sc_hd__xnor2_1 _15342_ (.A(_07985_),
    .B(_07986_),
    .Y(_07987_));
 sky130_fd_sc_hd__mux2_1 _15343_ (.A0(_07948_),
    .A1(_07987_),
    .S(_05335_),
    .X(_07988_));
 sky130_fd_sc_hd__nor2_1 _15344_ (.A(_05632_),
    .B(_07988_),
    .Y(_00477_));
 sky130_fd_sc_hd__or2b_1 _15345_ (.A(_07963_),
    .B_N(_07962_),
    .X(_07989_));
 sky130_fd_sc_hd__nand2_2 _15346_ (.A(_07624_),
    .B(_07637_),
    .Y(_07990_));
 sky130_fd_sc_hd__nor2_1 _15347_ (.A(_07619_),
    .B(_07824_),
    .Y(_07991_));
 sky130_fd_sc_hd__and3_1 _15348_ (.A(_07621_),
    .B(_07640_),
    .C(_07991_),
    .X(_07992_));
 sky130_fd_sc_hd__a21oi_1 _15349_ (.A1(_07621_),
    .A2(_07640_),
    .B1(_07991_),
    .Y(_07993_));
 sky130_fd_sc_hd__or2_1 _15350_ (.A(_07992_),
    .B(_07993_),
    .X(_07994_));
 sky130_fd_sc_hd__xor2_1 _15351_ (.A(_07990_),
    .B(_07994_),
    .X(_07995_));
 sky130_fd_sc_hd__a31o_1 _15352_ (.A1(_07622_),
    .A2(_07637_),
    .A3(_07959_),
    .B1(_07958_),
    .X(_07996_));
 sky130_fd_sc_hd__xor2_1 _15353_ (.A(_07995_),
    .B(_07996_),
    .X(_07997_));
 sky130_fd_sc_hd__nand2_1 _15354_ (.A(_07956_),
    .B(_07997_),
    .Y(_07998_));
 sky130_fd_sc_hd__or2_1 _15355_ (.A(_07956_),
    .B(_07997_),
    .X(_07999_));
 sky130_fd_sc_hd__nand2_1 _15356_ (.A(_07998_),
    .B(_07999_),
    .Y(_08000_));
 sky130_fd_sc_hd__a21o_1 _15357_ (.A1(_07989_),
    .A2(_07965_),
    .B1(_08000_),
    .X(_08001_));
 sky130_fd_sc_hd__nand3_1 _15358_ (.A(_07989_),
    .B(_07965_),
    .C(_08000_),
    .Y(_08002_));
 sky130_fd_sc_hd__nand2_1 _15359_ (.A(_08001_),
    .B(_08002_),
    .Y(_08003_));
 sky130_fd_sc_hd__a21o_1 _15360_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[11] ),
    .A2(_07924_),
    .B1(_07844_),
    .X(_08004_));
 sky130_fd_sc_hd__o21ba_2 _15361_ (.A1(_07881_),
    .A2(_07954_),
    .B1_N(_07916_),
    .X(_08005_));
 sky130_fd_sc_hd__xnor2_1 _15362_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[12] ),
    .B(_07845_),
    .Y(_08006_));
 sky130_fd_sc_hd__nor2_1 _15363_ (.A(_08005_),
    .B(_08006_),
    .Y(_08007_));
 sky130_fd_sc_hd__and2_1 _15364_ (.A(_08005_),
    .B(_08006_),
    .X(_08008_));
 sky130_fd_sc_hd__nor2_1 _15365_ (.A(_08007_),
    .B(_08008_),
    .Y(_08009_));
 sky130_fd_sc_hd__xnor2_1 _15366_ (.A(_08004_),
    .B(_08009_),
    .Y(_08010_));
 sky130_fd_sc_hd__xor2_1 _15367_ (.A(_08003_),
    .B(_08010_),
    .X(_08011_));
 sky130_fd_sc_hd__a21o_1 _15368_ (.A1(_07969_),
    .A2(_07975_),
    .B1(_07968_),
    .X(_08012_));
 sky130_fd_sc_hd__xnor2_1 _15369_ (.A(_08011_),
    .B(_08012_),
    .Y(_08013_));
 sky130_fd_sc_hd__or2b_1 _15370_ (.A(_07973_),
    .B_N(_07972_),
    .X(_08014_));
 sky130_fd_sc_hd__a21bo_1 _15371_ (.A1(_07971_),
    .A2(_07974_),
    .B1_N(_08014_),
    .X(_08015_));
 sky130_fd_sc_hd__xnor2_1 _15372_ (.A(_08013_),
    .B(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__or2b_1 _15373_ (.A(_07978_),
    .B_N(_07980_),
    .X(_08017_));
 sky130_fd_sc_hd__a21bo_1 _15374_ (.A1(_07976_),
    .A2(_07977_),
    .B1_N(_08017_),
    .X(_08018_));
 sky130_fd_sc_hd__and2_1 _15375_ (.A(_08016_),
    .B(_08018_),
    .X(_08019_));
 sky130_fd_sc_hd__nor2_1 _15376_ (.A(_08016_),
    .B(_08018_),
    .Y(_08020_));
 sky130_fd_sc_hd__nor2_1 _15377_ (.A(_08019_),
    .B(_08020_),
    .Y(_08021_));
 sky130_fd_sc_hd__xor2_2 _15378_ (.A(_07982_),
    .B(_08021_),
    .X(_08022_));
 sky130_fd_sc_hd__nand2_1 _15379_ (.A(_07949_),
    .B(_07984_),
    .Y(_08023_));
 sky130_fd_sc_hd__o21a_1 _15380_ (.A1(_07985_),
    .A2(_07986_),
    .B1(_08023_),
    .X(_08024_));
 sky130_fd_sc_hd__nor2_1 _15381_ (.A(_08022_),
    .B(_08024_),
    .Y(_08025_));
 sky130_fd_sc_hd__a21o_1 _15382_ (.A1(_08022_),
    .A2(_08024_),
    .B1(_06404_),
    .X(_08026_));
 sky130_fd_sc_hd__a2bb2o_1 _15383_ (.A1_N(_08025_),
    .A2_N(_08026_),
    .B1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[12] ),
    .B2(_07816_),
    .X(_08027_));
 sky130_fd_sc_hd__and2_1 _15384_ (.A(_07117_),
    .B(_08027_),
    .X(_08028_));
 sky130_fd_sc_hd__clkbuf_1 _15385_ (.A(_08028_),
    .X(_00478_));
 sky130_fd_sc_hd__nand2_1 _15386_ (.A(net974),
    .B(_05403_),
    .Y(_08029_));
 sky130_fd_sc_hd__nand2_1 _15387_ (.A(_07995_),
    .B(_07996_),
    .Y(_08030_));
 sky130_fd_sc_hd__nand2_1 _15388_ (.A(_07624_),
    .B(_07640_),
    .Y(_08031_));
 sky130_fd_sc_hd__o21a_1 _15389_ (.A1(_07622_),
    .A2(_07824_),
    .B1(_08031_),
    .X(_08032_));
 sky130_fd_sc_hd__nor3_1 _15390_ (.A(_07622_),
    .B(_07824_),
    .C(_08031_),
    .Y(_08033_));
 sky130_fd_sc_hd__nor2_1 _15391_ (.A(_08032_),
    .B(_08033_),
    .Y(_08034_));
 sky130_fd_sc_hd__xnor2_1 _15392_ (.A(_07990_),
    .B(_08034_),
    .Y(_08035_));
 sky130_fd_sc_hd__o21ba_1 _15393_ (.A1(_07990_),
    .A2(_07993_),
    .B1_N(_07992_),
    .X(_08036_));
 sky130_fd_sc_hd__xnor2_1 _15394_ (.A(_08035_),
    .B(_08036_),
    .Y(_08037_));
 sky130_fd_sc_hd__nand2_1 _15395_ (.A(_07956_),
    .B(_08037_),
    .Y(_08038_));
 sky130_fd_sc_hd__or2_1 _15396_ (.A(_07956_),
    .B(_08037_),
    .X(_08039_));
 sky130_fd_sc_hd__nand2_1 _15397_ (.A(_08038_),
    .B(_08039_),
    .Y(_08040_));
 sky130_fd_sc_hd__a21o_1 _15398_ (.A1(_08030_),
    .A2(_07998_),
    .B1(_08040_),
    .X(_08041_));
 sky130_fd_sc_hd__nand3_1 _15399_ (.A(_08030_),
    .B(_07998_),
    .C(_08040_),
    .Y(_08042_));
 sky130_fd_sc_hd__a21o_1 _15400_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[12] ),
    .A2(_07924_),
    .B1(_07844_),
    .X(_08043_));
 sky130_fd_sc_hd__xnor2_1 _15401_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[13] ),
    .B(_07924_),
    .Y(_08044_));
 sky130_fd_sc_hd__nor2_1 _15402_ (.A(_08005_),
    .B(_08044_),
    .Y(_08045_));
 sky130_fd_sc_hd__and2_1 _15403_ (.A(_08005_),
    .B(_08044_),
    .X(_08046_));
 sky130_fd_sc_hd__nor2_1 _15404_ (.A(_08045_),
    .B(_08046_),
    .Y(_08047_));
 sky130_fd_sc_hd__xor2_1 _15405_ (.A(_08043_),
    .B(_08047_),
    .X(_08048_));
 sky130_fd_sc_hd__and3_1 _15406_ (.A(_08041_),
    .B(_08042_),
    .C(_08048_),
    .X(_08049_));
 sky130_fd_sc_hd__a21oi_1 _15407_ (.A1(_08041_),
    .A2(_08042_),
    .B1(_08048_),
    .Y(_08050_));
 sky130_fd_sc_hd__nor2_1 _15408_ (.A(_08049_),
    .B(_08050_),
    .Y(_08051_));
 sky130_fd_sc_hd__o21ai_2 _15409_ (.A1(_08003_),
    .A2(_08010_),
    .B1(_08001_),
    .Y(_08052_));
 sky130_fd_sc_hd__xnor2_1 _15410_ (.A(_08051_),
    .B(_08052_),
    .Y(_08053_));
 sky130_fd_sc_hd__a21o_1 _15411_ (.A1(_08004_),
    .A2(_08009_),
    .B1(_08007_),
    .X(_08054_));
 sky130_fd_sc_hd__xnor2_1 _15412_ (.A(_08053_),
    .B(_08054_),
    .Y(_08055_));
 sky130_fd_sc_hd__or2b_1 _15413_ (.A(_08013_),
    .B_N(_08015_),
    .X(_08056_));
 sky130_fd_sc_hd__a21bo_1 _15414_ (.A1(_08011_),
    .A2(_08012_),
    .B1_N(_08056_),
    .X(_08057_));
 sky130_fd_sc_hd__nand2_1 _15415_ (.A(_08055_),
    .B(_08057_),
    .Y(_08058_));
 sky130_fd_sc_hd__or2_1 _15416_ (.A(_08055_),
    .B(_08057_),
    .X(_08059_));
 sky130_fd_sc_hd__and2_1 _15417_ (.A(_08058_),
    .B(_08059_),
    .X(_08060_));
 sky130_fd_sc_hd__xor2_2 _15418_ (.A(_08019_),
    .B(_08060_),
    .X(_08061_));
 sky130_fd_sc_hd__and2b_1 _15419_ (.A_N(_07982_),
    .B(_08021_),
    .X(_08062_));
 sky130_fd_sc_hd__o21bai_2 _15420_ (.A1(_08022_),
    .A2(_08024_),
    .B1_N(_08062_),
    .Y(_08063_));
 sky130_fd_sc_hd__a21oi_1 _15421_ (.A1(_08061_),
    .A2(_08063_),
    .B1(_06734_),
    .Y(_08064_));
 sky130_fd_sc_hd__o21ai_1 _15422_ (.A1(_08061_),
    .A2(_08063_),
    .B1(_08064_),
    .Y(_08065_));
 sky130_fd_sc_hd__a21oi_1 _15423_ (.A1(_08029_),
    .A2(_08065_),
    .B1(_05440_),
    .Y(_00479_));
 sky130_fd_sc_hd__buf_4 _15424_ (.A(_05353_),
    .X(_08066_));
 sky130_fd_sc_hd__a21oi_1 _15425_ (.A1(_08030_),
    .A2(_07998_),
    .B1(_08040_),
    .Y(_08067_));
 sky130_fd_sc_hd__or2b_1 _15426_ (.A(_08036_),
    .B_N(_08035_),
    .X(_08068_));
 sky130_fd_sc_hd__and3_1 _15427_ (.A(_07624_),
    .B(_07640_),
    .C(_07637_),
    .X(_08069_));
 sky130_fd_sc_hd__o21ba_1 _15428_ (.A1(_07990_),
    .A2(_08032_),
    .B1_N(_08033_),
    .X(_08070_));
 sky130_fd_sc_hd__o21a_1 _15429_ (.A1(_07624_),
    .A2(_07824_),
    .B1(_08031_),
    .X(_08071_));
 sky130_fd_sc_hd__a2bb2o_1 _15430_ (.A1_N(_08069_),
    .A2_N(_08070_),
    .B1(_07990_),
    .B2(_08071_),
    .X(_08072_));
 sky130_fd_sc_hd__xor2_1 _15431_ (.A(_07956_),
    .B(_08072_),
    .X(_08073_));
 sky130_fd_sc_hd__a21oi_1 _15432_ (.A1(_08068_),
    .A2(_08038_),
    .B1(_08073_),
    .Y(_08074_));
 sky130_fd_sc_hd__nand3_1 _15433_ (.A(_08068_),
    .B(_08038_),
    .C(_08073_),
    .Y(_08075_));
 sky130_fd_sc_hd__or2b_1 _15434_ (.A(_08074_),
    .B_N(_08075_),
    .X(_08076_));
 sky130_fd_sc_hd__a21oi_1 _15435_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[13] ),
    .A2(_07924_),
    .B1(_07844_),
    .Y(_08077_));
 sky130_fd_sc_hd__xnor2_1 _15436_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[14] ),
    .B(_07924_),
    .Y(_08078_));
 sky130_fd_sc_hd__nor2_1 _15437_ (.A(_08005_),
    .B(_08078_),
    .Y(_08079_));
 sky130_fd_sc_hd__and2_1 _15438_ (.A(_08005_),
    .B(_08078_),
    .X(_08080_));
 sky130_fd_sc_hd__nor2_1 _15439_ (.A(_08079_),
    .B(_08080_),
    .Y(_08081_));
 sky130_fd_sc_hd__xnor2_1 _15440_ (.A(_08077_),
    .B(_08081_),
    .Y(_08082_));
 sky130_fd_sc_hd__xnor2_1 _15441_ (.A(_08076_),
    .B(_08082_),
    .Y(_08083_));
 sky130_fd_sc_hd__o21ai_1 _15442_ (.A1(_08067_),
    .A2(_08049_),
    .B1(_08083_),
    .Y(_08084_));
 sky130_fd_sc_hd__or3_1 _15443_ (.A(_08067_),
    .B(_08049_),
    .C(_08083_),
    .X(_08085_));
 sky130_fd_sc_hd__nand2_1 _15444_ (.A(_08084_),
    .B(_08085_),
    .Y(_08086_));
 sky130_fd_sc_hd__a21oi_2 _15445_ (.A1(_08043_),
    .A2(_08047_),
    .B1(_08045_),
    .Y(_08087_));
 sky130_fd_sc_hd__xnor2_2 _15446_ (.A(_08086_),
    .B(_08087_),
    .Y(_08088_));
 sky130_fd_sc_hd__or2b_1 _15447_ (.A(_08053_),
    .B_N(_08054_),
    .X(_08089_));
 sky130_fd_sc_hd__a21boi_2 _15448_ (.A1(_08051_),
    .A2(_08052_),
    .B1_N(_08089_),
    .Y(_08090_));
 sky130_fd_sc_hd__xnor2_1 _15449_ (.A(_08088_),
    .B(_08090_),
    .Y(_08091_));
 sky130_fd_sc_hd__nor2_1 _15450_ (.A(_08058_),
    .B(_08091_),
    .Y(_08092_));
 sky130_fd_sc_hd__and2_1 _15451_ (.A(_08058_),
    .B(_08091_),
    .X(_08093_));
 sky130_fd_sc_hd__nor2_1 _15452_ (.A(_08092_),
    .B(_08093_),
    .Y(_08094_));
 sky130_fd_sc_hd__a32o_1 _15453_ (.A1(_08016_),
    .A2(_08018_),
    .A3(_08060_),
    .B1(_08061_),
    .B2(_08063_),
    .X(_08095_));
 sky130_fd_sc_hd__nand2_1 _15454_ (.A(_08094_),
    .B(_08095_),
    .Y(_08096_));
 sky130_fd_sc_hd__o21a_1 _15455_ (.A1(_08094_),
    .A2(_08095_),
    .B1(_05315_),
    .X(_08097_));
 sky130_fd_sc_hd__a22o_1 _15456_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[14] ),
    .A2(_08066_),
    .B1(_08096_),
    .B2(_08097_),
    .X(_08098_));
 sky130_fd_sc_hd__and2_1 _15457_ (.A(_07117_),
    .B(_08098_),
    .X(_08099_));
 sky130_fd_sc_hd__clkbuf_1 _15458_ (.A(_08099_),
    .X(_00480_));
 sky130_fd_sc_hd__and2_1 _15459_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[15] ),
    .B(_07576_),
    .X(_08100_));
 sky130_fd_sc_hd__a21oi_1 _15460_ (.A1(_08075_),
    .A2(_08082_),
    .B1(_08074_),
    .Y(_08101_));
 sky130_fd_sc_hd__and2b_1 _15461_ (.A_N(_07956_),
    .B(_08072_),
    .X(_08102_));
 sky130_fd_sc_hd__a21o_1 _15462_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[14] ),
    .A2(_07924_),
    .B1(_07844_),
    .X(_08103_));
 sky130_fd_sc_hd__xnor2_2 _15463_ (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[15] ),
    .B(_07924_),
    .Y(_08104_));
 sky130_fd_sc_hd__xnor2_1 _15464_ (.A(_08005_),
    .B(_08104_),
    .Y(_08105_));
 sky130_fd_sc_hd__xnor2_1 _15465_ (.A(_08103_),
    .B(_08105_),
    .Y(_08106_));
 sky130_fd_sc_hd__or2_1 _15466_ (.A(_08102_),
    .B(_08106_),
    .X(_08107_));
 sky130_fd_sc_hd__nand2_1 _15467_ (.A(_08102_),
    .B(_08106_),
    .Y(_08108_));
 sky130_fd_sc_hd__and2_1 _15468_ (.A(_08107_),
    .B(_08108_),
    .X(_08109_));
 sky130_fd_sc_hd__xnor2_1 _15469_ (.A(_08101_),
    .B(_08109_),
    .Y(_08110_));
 sky130_fd_sc_hd__o21ba_1 _15470_ (.A1(_08077_),
    .A2(_08080_),
    .B1_N(_08079_),
    .X(_08111_));
 sky130_fd_sc_hd__xnor2_1 _15471_ (.A(_08110_),
    .B(_08111_),
    .Y(_08112_));
 sky130_fd_sc_hd__o21a_1 _15472_ (.A1(_08086_),
    .A2(_08087_),
    .B1(_08084_),
    .X(_08113_));
 sky130_fd_sc_hd__or2_1 _15473_ (.A(_08112_),
    .B(_08113_),
    .X(_08114_));
 sky130_fd_sc_hd__nand2_1 _15474_ (.A(_08112_),
    .B(_08113_),
    .Y(_08115_));
 sky130_fd_sc_hd__and4bb_1 _15475_ (.A_N(_08088_),
    .B_N(_08090_),
    .C(_08114_),
    .D(_08115_),
    .X(_08116_));
 sky130_fd_sc_hd__and2_1 _15476_ (.A(_08114_),
    .B(_08115_),
    .X(_08117_));
 sky130_fd_sc_hd__o21ba_1 _15477_ (.A1(_08088_),
    .A2(_08090_),
    .B1_N(_08117_),
    .X(_08118_));
 sky130_fd_sc_hd__a21oi_1 _15478_ (.A1(_08094_),
    .A2(_08095_),
    .B1(_08092_),
    .Y(_08119_));
 sky130_fd_sc_hd__nor2_1 _15479_ (.A(_08116_),
    .B(_08118_),
    .Y(_08120_));
 sky130_fd_sc_hd__a211o_1 _15480_ (.A1(_08094_),
    .A2(_08095_),
    .B1(_08120_),
    .C1(_08092_),
    .X(_08121_));
 sky130_fd_sc_hd__o311a_1 _15481_ (.A1(_08116_),
    .A2(_08118_),
    .A3(_08119_),
    .B1(_08121_),
    .C1(_05313_),
    .X(_08122_));
 sky130_fd_sc_hd__o21a_1 _15482_ (.A1(_08100_),
    .A2(_08122_),
    .B1(_04870_),
    .X(_00481_));
 sky130_fd_sc_hd__or2_1 _15483_ (.A(_08101_),
    .B(_08109_),
    .X(_08123_));
 sky130_fd_sc_hd__o21a_1 _15484_ (.A1(_08110_),
    .A2(_08111_),
    .B1(_08123_),
    .X(_08124_));
 sky130_fd_sc_hd__xnor2_1 _15485_ (.A(_08107_),
    .B(_08124_),
    .Y(_08125_));
 sky130_fd_sc_hd__a21o_1 _15486_ (.A1(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[15] ),
    .A2(_07924_),
    .B1(_07844_),
    .X(_08126_));
 sky130_fd_sc_hd__o21a_1 _15487_ (.A1(_08005_),
    .A2(_08104_),
    .B1(_08103_),
    .X(_08127_));
 sky130_fd_sc_hd__a21oi_1 _15488_ (.A1(_08005_),
    .A2(_08104_),
    .B1(_08127_),
    .Y(_08128_));
 sky130_fd_sc_hd__xnor2_1 _15489_ (.A(_08114_),
    .B(_08128_),
    .Y(_08129_));
 sky130_fd_sc_hd__xnor2_1 _15490_ (.A(_08126_),
    .B(_08129_),
    .Y(_08130_));
 sky130_fd_sc_hd__xnor2_1 _15491_ (.A(_08125_),
    .B(_08130_),
    .Y(_08131_));
 sky130_fd_sc_hd__nor2_1 _15492_ (.A(_08116_),
    .B(_08131_),
    .Y(_08132_));
 sky130_fd_sc_hd__o31a_1 _15493_ (.A1(_08116_),
    .A2(_08118_),
    .A3(_08119_),
    .B1(_08132_),
    .X(_08133_));
 sky130_fd_sc_hd__or2_1 _15494_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[16] ),
    .B(_07866_),
    .X(_08134_));
 sky130_fd_sc_hd__o211a_1 _15495_ (.A1(_06848_),
    .A2(_08133_),
    .B1(_08134_),
    .C1(_07643_),
    .X(_00482_));
 sky130_fd_sc_hd__clkbuf_4 _15496_ (.A(\top_inst.grid_inst.data_path_wires[7][0] ),
    .X(_08135_));
 sky130_fd_sc_hd__or2_1 _15497_ (.A(_08135_),
    .B(_06620_),
    .X(_08136_));
 sky130_fd_sc_hd__o211a_1 _15498_ (.A1(_07606_),
    .A2(_06634_),
    .B1(_08136_),
    .C1(_07643_),
    .X(_00483_));
 sky130_fd_sc_hd__buf_4 _15499_ (.A(\top_inst.grid_inst.data_path_wires[7][1] ),
    .X(_08137_));
 sky130_fd_sc_hd__or2_1 _15500_ (.A(_08137_),
    .B(_06620_),
    .X(_08138_));
 sky130_fd_sc_hd__o211a_1 _15501_ (.A1(_07608_),
    .A2(_06634_),
    .B1(_08138_),
    .C1(_07643_),
    .X(_00484_));
 sky130_fd_sc_hd__clkbuf_4 _15502_ (.A(\top_inst.grid_inst.data_path_wires[7][2] ),
    .X(_08139_));
 sky130_fd_sc_hd__buf_2 _15503_ (.A(_06619_),
    .X(_08140_));
 sky130_fd_sc_hd__or2_1 _15504_ (.A(_08139_),
    .B(_08140_),
    .X(_08141_));
 sky130_fd_sc_hd__clkbuf_4 _15505_ (.A(_07617_),
    .X(_08142_));
 sky130_fd_sc_hd__o211a_1 _15506_ (.A1(_07610_),
    .A2(_06634_),
    .B1(_08141_),
    .C1(_08142_),
    .X(_00485_));
 sky130_fd_sc_hd__buf_4 _15507_ (.A(\top_inst.grid_inst.data_path_wires[7][3] ),
    .X(_08143_));
 sky130_fd_sc_hd__or2_1 _15508_ (.A(_08143_),
    .B(_08140_),
    .X(_08144_));
 sky130_fd_sc_hd__o211a_1 _15509_ (.A1(_07613_),
    .A2(_06634_),
    .B1(_08144_),
    .C1(_08142_),
    .X(_00486_));
 sky130_fd_sc_hd__inv_2 _15510_ (.A(\top_inst.grid_inst.data_path_wires[7][4] ),
    .Y(_08145_));
 sky130_fd_sc_hd__nand2_1 _15511_ (.A(_08145_),
    .B(_04859_),
    .Y(_08146_));
 sky130_fd_sc_hd__o211a_1 _15512_ (.A1(_07615_),
    .A2(_06634_),
    .B1(_08146_),
    .C1(_08142_),
    .X(_00487_));
 sky130_fd_sc_hd__buf_4 _15513_ (.A(\top_inst.grid_inst.data_path_wires[7][5] ),
    .X(_08147_));
 sky130_fd_sc_hd__or2_1 _15514_ (.A(_08147_),
    .B(_08140_),
    .X(_08148_));
 sky130_fd_sc_hd__o211a_1 _15515_ (.A1(_07619_),
    .A2(_06634_),
    .B1(_08148_),
    .C1(_08142_),
    .X(_00488_));
 sky130_fd_sc_hd__buf_2 _15516_ (.A(\top_inst.grid_inst.data_path_wires[7][6] ),
    .X(_08149_));
 sky130_fd_sc_hd__buf_4 _15517_ (.A(_08149_),
    .X(_08150_));
 sky130_fd_sc_hd__or2_1 _15518_ (.A(_08150_),
    .B(_08140_),
    .X(_08151_));
 sky130_fd_sc_hd__o211a_1 _15519_ (.A1(_07622_),
    .A2(_06634_),
    .B1(_08151_),
    .C1(_08142_),
    .X(_00489_));
 sky130_fd_sc_hd__buf_4 _15520_ (.A(\top_inst.grid_inst.data_path_wires[7][7] ),
    .X(_08152_));
 sky130_fd_sc_hd__or2_1 _15521_ (.A(_08152_),
    .B(_08140_),
    .X(_08153_));
 sky130_fd_sc_hd__o211a_1 _15522_ (.A1(_07624_),
    .A2(_06634_),
    .B1(_08153_),
    .C1(_08142_),
    .X(_00490_));
 sky130_fd_sc_hd__buf_2 _15523_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[0] ),
    .X(_08154_));
 sky130_fd_sc_hd__clkbuf_4 _15524_ (.A(_08154_),
    .X(_08155_));
 sky130_fd_sc_hd__or2_1 _15525_ (.A(_08155_),
    .B(_07641_),
    .X(_08156_));
 sky130_fd_sc_hd__o211a_1 _15526_ (.A1(_08135_),
    .A2(_07639_),
    .B1(_08156_),
    .C1(_08142_),
    .X(_00491_));
 sky130_fd_sc_hd__clkbuf_4 _15527_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[1] ),
    .X(_08157_));
 sky130_fd_sc_hd__or2_1 _15528_ (.A(_08157_),
    .B(_07641_),
    .X(_08158_));
 sky130_fd_sc_hd__o211a_1 _15529_ (.A1(_08137_),
    .A2(_07639_),
    .B1(_08158_),
    .C1(_08142_),
    .X(_00492_));
 sky130_fd_sc_hd__buf_4 _15530_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[2] ),
    .X(_08159_));
 sky130_fd_sc_hd__or2_1 _15531_ (.A(_08159_),
    .B(_07641_),
    .X(_08160_));
 sky130_fd_sc_hd__o211a_1 _15532_ (.A1(_08139_),
    .A2(_07639_),
    .B1(_08160_),
    .C1(_08142_),
    .X(_00493_));
 sky130_fd_sc_hd__clkbuf_4 _15533_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[3] ),
    .X(_08161_));
 sky130_fd_sc_hd__or2_1 _15534_ (.A(_08161_),
    .B(_07641_),
    .X(_08162_));
 sky130_fd_sc_hd__o211a_1 _15535_ (.A1(_08143_),
    .A2(_07639_),
    .B1(_08162_),
    .C1(_08142_),
    .X(_00494_));
 sky130_fd_sc_hd__buf_4 _15536_ (.A(\top_inst.grid_inst.data_path_wires[7][4] ),
    .X(_08163_));
 sky130_fd_sc_hd__clkbuf_4 _15537_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[4] ),
    .X(_08164_));
 sky130_fd_sc_hd__or2_1 _15538_ (.A(_08164_),
    .B(_07641_),
    .X(_08165_));
 sky130_fd_sc_hd__clkbuf_4 _15539_ (.A(_07617_),
    .X(_08166_));
 sky130_fd_sc_hd__o211a_1 _15540_ (.A1(_08163_),
    .A2(_07639_),
    .B1(_08165_),
    .C1(_08166_),
    .X(_00495_));
 sky130_fd_sc_hd__clkbuf_4 _15541_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[5] ),
    .X(_08167_));
 sky130_fd_sc_hd__or2_1 _15542_ (.A(_08167_),
    .B(_07641_),
    .X(_08168_));
 sky130_fd_sc_hd__o211a_1 _15543_ (.A1(_08147_),
    .A2(_07639_),
    .B1(_08168_),
    .C1(_08166_),
    .X(_00496_));
 sky130_fd_sc_hd__buf_2 _15544_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[6] ),
    .X(_08169_));
 sky130_fd_sc_hd__or2_1 _15545_ (.A(_08169_),
    .B(_07641_),
    .X(_08170_));
 sky130_fd_sc_hd__o211a_1 _15546_ (.A1(_08150_),
    .A2(_07639_),
    .B1(_08170_),
    .C1(_08166_),
    .X(_00497_));
 sky130_fd_sc_hd__or2_1 _15547_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[7] ),
    .B(_07641_),
    .X(_08171_));
 sky130_fd_sc_hd__o211a_1 _15548_ (.A1(_08152_),
    .A2(_07639_),
    .B1(_08171_),
    .C1(_08166_),
    .X(_00498_));
 sky130_fd_sc_hd__and3_1 _15549_ (.A(_08135_),
    .B(_08155_),
    .C(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[0] ),
    .X(_08172_));
 sky130_fd_sc_hd__a21oi_1 _15550_ (.A1(_08135_),
    .A2(_08155_),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[0] ),
    .Y(_08173_));
 sky130_fd_sc_hd__o21ai_1 _15551_ (.A1(_08172_),
    .A2(_08173_),
    .B1(_05336_),
    .Y(_08174_));
 sky130_fd_sc_hd__o211a_1 _15552_ (.A1(net1075),
    .A2(_06660_),
    .B1(_08174_),
    .C1(_08166_),
    .X(_00499_));
 sky130_fd_sc_hd__a22o_1 _15553_ (.A1(_08135_),
    .A2(_08157_),
    .B1(_08155_),
    .B2(_08137_),
    .X(_08175_));
 sky130_fd_sc_hd__nand4_2 _15554_ (.A(_08137_),
    .B(_08135_),
    .C(_08157_),
    .D(_08155_),
    .Y(_08176_));
 sky130_fd_sc_hd__nand3_1 _15555_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[1] ),
    .B(_08175_),
    .C(_08176_),
    .Y(_08177_));
 sky130_fd_sc_hd__a21o_1 _15556_ (.A1(_08175_),
    .A2(_08176_),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[1] ),
    .X(_08178_));
 sky130_fd_sc_hd__a21oi_1 _15557_ (.A1(_08177_),
    .A2(_08178_),
    .B1(_08172_),
    .Y(_08179_));
 sky130_fd_sc_hd__and3_1 _15558_ (.A(_08172_),
    .B(_08177_),
    .C(_08178_),
    .X(_08180_));
 sky130_fd_sc_hd__buf_6 _15559_ (.A(_05335_),
    .X(_08181_));
 sky130_fd_sc_hd__o21ai_1 _15560_ (.A1(_08179_),
    .A2(_08180_),
    .B1(_08181_),
    .Y(_08182_));
 sky130_fd_sc_hd__o211a_1 _15561_ (.A1(net1027),
    .A2(_06660_),
    .B1(_08182_),
    .C1(_08166_),
    .X(_00500_));
 sky130_fd_sc_hd__buf_8 _15562_ (.A(_05787_),
    .X(_08183_));
 sky130_fd_sc_hd__a22o_1 _15563_ (.A1(_08137_),
    .A2(_08157_),
    .B1(_08155_),
    .B2(_08139_),
    .X(_08184_));
 sky130_fd_sc_hd__nand4_1 _15564_ (.A(_08139_),
    .B(_08137_),
    .C(_08157_),
    .D(_08155_),
    .Y(_08185_));
 sky130_fd_sc_hd__nand2_1 _15565_ (.A(_08184_),
    .B(_08185_),
    .Y(_08186_));
 sky130_fd_sc_hd__xor2_1 _15566_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[2] ),
    .B(_08186_),
    .X(_08187_));
 sky130_fd_sc_hd__nand2_1 _15567_ (.A(_08176_),
    .B(_08177_),
    .Y(_08188_));
 sky130_fd_sc_hd__xnor2_1 _15568_ (.A(_08187_),
    .B(_08188_),
    .Y(_08189_));
 sky130_fd_sc_hd__and2_1 _15569_ (.A(_08135_),
    .B(_08159_),
    .X(_08190_));
 sky130_fd_sc_hd__or2_1 _15570_ (.A(_08189_),
    .B(_08190_),
    .X(_08191_));
 sky130_fd_sc_hd__nand2_1 _15571_ (.A(_08189_),
    .B(_08190_),
    .Y(_08192_));
 sky130_fd_sc_hd__and2_1 _15572_ (.A(_08191_),
    .B(_08192_),
    .X(_08193_));
 sky130_fd_sc_hd__or2_1 _15573_ (.A(_08180_),
    .B(_08193_),
    .X(_08194_));
 sky130_fd_sc_hd__nand2_1 _15574_ (.A(_08180_),
    .B(_08193_),
    .Y(_08195_));
 sky130_fd_sc_hd__a21o_1 _15575_ (.A1(_08194_),
    .A2(_08195_),
    .B1(_06682_),
    .X(_08196_));
 sky130_fd_sc_hd__o211a_1 _15576_ (.A1(net1079),
    .A2(_08183_),
    .B1(_08196_),
    .C1(_08166_),
    .X(_00501_));
 sky130_fd_sc_hd__clkbuf_4 _15577_ (.A(_04869_),
    .X(_08197_));
 sky130_fd_sc_hd__or2b_1 _15578_ (.A(_08187_),
    .B_N(_08188_),
    .X(_08198_));
 sky130_fd_sc_hd__a22o_1 _15579_ (.A1(_08135_),
    .A2(_08161_),
    .B1(_08159_),
    .B2(_08137_),
    .X(_08199_));
 sky130_fd_sc_hd__and3_1 _15580_ (.A(\top_inst.grid_inst.data_path_wires[7][1] ),
    .B(\top_inst.grid_inst.data_path_wires[7][0] ),
    .C(_08161_),
    .X(_08200_));
 sky130_fd_sc_hd__nand2_2 _15581_ (.A(_08159_),
    .B(_08200_),
    .Y(_08201_));
 sky130_fd_sc_hd__nand2_1 _15582_ (.A(_08199_),
    .B(_08201_),
    .Y(_08202_));
 sky130_fd_sc_hd__a22o_1 _15583_ (.A1(_08139_),
    .A2(_08157_),
    .B1(_08155_),
    .B2(_08143_),
    .X(_08203_));
 sky130_fd_sc_hd__nand4_1 _15584_ (.A(_08143_),
    .B(_08139_),
    .C(_08157_),
    .D(_08155_),
    .Y(_08204_));
 sky130_fd_sc_hd__and3_1 _15585_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[3] ),
    .B(_08203_),
    .C(_08204_),
    .X(_08205_));
 sky130_fd_sc_hd__a21oi_1 _15586_ (.A1(_08203_),
    .A2(_08204_),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[3] ),
    .Y(_08206_));
 sky130_fd_sc_hd__or2_1 _15587_ (.A(_08205_),
    .B(_08206_),
    .X(_08207_));
 sky130_fd_sc_hd__a21boi_2 _15588_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[2] ),
    .A2(_08184_),
    .B1_N(_08185_),
    .Y(_08208_));
 sky130_fd_sc_hd__xnor2_1 _15589_ (.A(_08207_),
    .B(_08208_),
    .Y(_08209_));
 sky130_fd_sc_hd__xnor2_1 _15590_ (.A(_08202_),
    .B(_08209_),
    .Y(_08210_));
 sky130_fd_sc_hd__a21o_1 _15591_ (.A1(_08198_),
    .A2(_08192_),
    .B1(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__inv_2 _15592_ (.A(_08211_),
    .Y(_08212_));
 sky130_fd_sc_hd__and3_1 _15593_ (.A(_08198_),
    .B(_08192_),
    .C(_08210_),
    .X(_08213_));
 sky130_fd_sc_hd__or3_1 _15594_ (.A(_08195_),
    .B(_08212_),
    .C(_08213_),
    .X(_08214_));
 sky130_fd_sc_hd__o21ai_1 _15595_ (.A1(_08212_),
    .A2(_08213_),
    .B1(_08195_),
    .Y(_08215_));
 sky130_fd_sc_hd__and2_1 _15596_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[3] ),
    .B(_05326_),
    .X(_08216_));
 sky130_fd_sc_hd__a31o_1 _15597_ (.A1(_05887_),
    .A2(_08214_),
    .A3(_08215_),
    .B1(_08216_),
    .X(_08217_));
 sky130_fd_sc_hd__and2_1 _15598_ (.A(_08197_),
    .B(_08217_),
    .X(_08218_));
 sky130_fd_sc_hd__clkbuf_1 _15599_ (.A(_08218_),
    .X(_00502_));
 sky130_fd_sc_hd__a22o_1 _15600_ (.A1(\top_inst.grid_inst.data_path_wires[7][3] ),
    .A2(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[1] ),
    .B1(_08154_),
    .B2(\top_inst.grid_inst.data_path_wires[7][4] ),
    .X(_08219_));
 sky130_fd_sc_hd__nand4_1 _15601_ (.A(_08163_),
    .B(\top_inst.grid_inst.data_path_wires[7][3] ),
    .C(_08157_),
    .D(_08154_),
    .Y(_08220_));
 sky130_fd_sc_hd__nand2_1 _15602_ (.A(_08219_),
    .B(_08220_),
    .Y(_08221_));
 sky130_fd_sc_hd__xor2_2 _15603_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[4] ),
    .B(_08221_),
    .X(_08222_));
 sky130_fd_sc_hd__xor2_2 _15604_ (.A(_08201_),
    .B(_08222_),
    .X(_08223_));
 sky130_fd_sc_hd__a21bo_1 _15605_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[3] ),
    .A2(_08203_),
    .B1_N(_08204_),
    .X(_08224_));
 sky130_fd_sc_hd__xnor2_2 _15606_ (.A(_08223_),
    .B(_08224_),
    .Y(_08225_));
 sky130_fd_sc_hd__nand2_1 _15607_ (.A(_08139_),
    .B(_08159_),
    .Y(_08226_));
 sky130_fd_sc_hd__a22o_1 _15608_ (.A1(\top_inst.grid_inst.data_path_wires[7][0] ),
    .A2(_08164_),
    .B1(_08161_),
    .B2(\top_inst.grid_inst.data_path_wires[7][1] ),
    .X(_08227_));
 sky130_fd_sc_hd__a21bo_1 _15609_ (.A1(_08164_),
    .A2(_08200_),
    .B1_N(_08227_),
    .X(_08228_));
 sky130_fd_sc_hd__xor2_2 _15610_ (.A(_08226_),
    .B(_08228_),
    .X(_08229_));
 sky130_fd_sc_hd__xor2_2 _15611_ (.A(_08225_),
    .B(_08229_),
    .X(_08230_));
 sky130_fd_sc_hd__or2_1 _15612_ (.A(_08202_),
    .B(_08209_),
    .X(_08231_));
 sky130_fd_sc_hd__o21ai_2 _15613_ (.A1(_08207_),
    .A2(_08208_),
    .B1(_08231_),
    .Y(_08232_));
 sky130_fd_sc_hd__xor2_2 _15614_ (.A(_08230_),
    .B(_08232_),
    .X(_08233_));
 sky130_fd_sc_hd__nand2_1 _15615_ (.A(_08211_),
    .B(_08214_),
    .Y(_08234_));
 sky130_fd_sc_hd__nor2_1 _15616_ (.A(_08233_),
    .B(_08234_),
    .Y(_08235_));
 sky130_fd_sc_hd__a21o_1 _15617_ (.A1(_08233_),
    .A2(_08234_),
    .B1(_07057_),
    .X(_08236_));
 sky130_fd_sc_hd__o221a_1 _15618_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[4] ),
    .A2(_07048_),
    .B1(_08235_),
    .B2(_08236_),
    .C1(_07708_),
    .X(_00503_));
 sky130_fd_sc_hd__nor2_1 _15619_ (.A(_08214_),
    .B(_08233_),
    .Y(_08237_));
 sky130_fd_sc_hd__and2b_1 _15620_ (.A_N(_08225_),
    .B(_08229_),
    .X(_08238_));
 sky130_fd_sc_hd__nand2_1 _15621_ (.A(_08135_),
    .B(_08167_),
    .Y(_08239_));
 sky130_fd_sc_hd__a22o_1 _15622_ (.A1(\top_inst.grid_inst.data_path_wires[7][1] ),
    .A2(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[7][2] ),
    .X(_08240_));
 sky130_fd_sc_hd__nand4_4 _15623_ (.A(\top_inst.grid_inst.data_path_wires[7][2] ),
    .B(\top_inst.grid_inst.data_path_wires[7][1] ),
    .C(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[3] ),
    .Y(_08241_));
 sky130_fd_sc_hd__a22o_1 _15624_ (.A1(_08143_),
    .A2(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[2] ),
    .B1(_08240_),
    .B2(_08241_),
    .X(_08242_));
 sky130_fd_sc_hd__nand4_2 _15625_ (.A(_08143_),
    .B(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[2] ),
    .C(_08240_),
    .D(_08241_),
    .Y(_08243_));
 sky130_fd_sc_hd__nand2_1 _15626_ (.A(_08242_),
    .B(_08243_),
    .Y(_08244_));
 sky130_fd_sc_hd__or2_1 _15627_ (.A(_08239_),
    .B(_08244_),
    .X(_08245_));
 sky130_fd_sc_hd__nand2_1 _15628_ (.A(_08239_),
    .B(_08244_),
    .Y(_08246_));
 sky130_fd_sc_hd__and2_1 _15629_ (.A(_08245_),
    .B(_08246_),
    .X(_08247_));
 sky130_fd_sc_hd__a21boi_2 _15630_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[4] ),
    .A2(_08219_),
    .B1_N(_08220_),
    .Y(_08248_));
 sky130_fd_sc_hd__a32o_1 _15631_ (.A1(_08139_),
    .A2(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[2] ),
    .A3(_08227_),
    .B1(_08200_),
    .B2(_08164_),
    .X(_08249_));
 sky130_fd_sc_hd__a22o_1 _15632_ (.A1(\top_inst.grid_inst.data_path_wires[7][4] ),
    .A2(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[1] ),
    .B1(_08154_),
    .B2(\top_inst.grid_inst.data_path_wires[7][5] ),
    .X(_08250_));
 sky130_fd_sc_hd__nand4_1 _15633_ (.A(\top_inst.grid_inst.data_path_wires[7][5] ),
    .B(\top_inst.grid_inst.data_path_wires[7][4] ),
    .C(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[1] ),
    .D(_08154_),
    .Y(_08251_));
 sky130_fd_sc_hd__nand2_1 _15634_ (.A(_08250_),
    .B(_08251_),
    .Y(_08252_));
 sky130_fd_sc_hd__xor2_2 _15635_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[5] ),
    .B(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__xnor2_2 _15636_ (.A(_08249_),
    .B(_08253_),
    .Y(_08254_));
 sky130_fd_sc_hd__xnor2_2 _15637_ (.A(_08248_),
    .B(_08254_),
    .Y(_08255_));
 sky130_fd_sc_hd__xor2_2 _15638_ (.A(_08247_),
    .B(_08255_),
    .X(_08256_));
 sky130_fd_sc_hd__xor2_2 _15639_ (.A(_08238_),
    .B(_08256_),
    .X(_08257_));
 sky130_fd_sc_hd__nor2_1 _15640_ (.A(_08201_),
    .B(_08222_),
    .Y(_08258_));
 sky130_fd_sc_hd__a21o_1 _15641_ (.A1(_08223_),
    .A2(_08224_),
    .B1(_08258_),
    .X(_08259_));
 sky130_fd_sc_hd__xnor2_2 _15642_ (.A(_08257_),
    .B(_08259_),
    .Y(_08260_));
 sky130_fd_sc_hd__or2b_1 _15643_ (.A(_08230_),
    .B_N(_08232_),
    .X(_08261_));
 sky130_fd_sc_hd__o21a_1 _15644_ (.A1(_08211_),
    .A2(_08233_),
    .B1(_08261_),
    .X(_08262_));
 sky130_fd_sc_hd__xor2_1 _15645_ (.A(_08260_),
    .B(_08262_),
    .X(_08263_));
 sky130_fd_sc_hd__nand2_1 _15646_ (.A(_08237_),
    .B(_08263_),
    .Y(_08264_));
 sky130_fd_sc_hd__buf_6 _15647_ (.A(_05311_),
    .X(_08265_));
 sky130_fd_sc_hd__o21a_1 _15648_ (.A1(_08237_),
    .A2(_08263_),
    .B1(_08265_),
    .X(_08266_));
 sky130_fd_sc_hd__a22o_1 _15649_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[5] ),
    .A2(_08066_),
    .B1(_08264_),
    .B2(_08266_),
    .X(_08267_));
 sky130_fd_sc_hd__and2_1 _15650_ (.A(_08197_),
    .B(_08267_),
    .X(_08268_));
 sky130_fd_sc_hd__clkbuf_1 _15651_ (.A(_08268_),
    .X(_00504_));
 sky130_fd_sc_hd__nor2_1 _15652_ (.A(_08261_),
    .B(_08260_),
    .Y(_08269_));
 sky130_fd_sc_hd__nand2_1 _15653_ (.A(_08238_),
    .B(_08256_),
    .Y(_08270_));
 sky130_fd_sc_hd__nand2_1 _15654_ (.A(_08257_),
    .B(_08259_),
    .Y(_08271_));
 sky130_fd_sc_hd__or2b_1 _15655_ (.A(_08253_),
    .B_N(_08249_),
    .X(_08272_));
 sky130_fd_sc_hd__or2b_1 _15656_ (.A(_08248_),
    .B_N(_08254_),
    .X(_08273_));
 sky130_fd_sc_hd__a22o_1 _15657_ (.A1(\top_inst.grid_inst.data_path_wires[7][0] ),
    .A2(_08169_),
    .B1(_08167_),
    .B2(_08137_),
    .X(_08274_));
 sky130_fd_sc_hd__nand4_2 _15658_ (.A(_08137_),
    .B(\top_inst.grid_inst.data_path_wires[7][0] ),
    .C(_08169_),
    .D(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[5] ),
    .Y(_08275_));
 sky130_fd_sc_hd__nand2_1 _15659_ (.A(_08274_),
    .B(_08275_),
    .Y(_08276_));
 sky130_fd_sc_hd__a22o_1 _15660_ (.A1(\top_inst.grid_inst.data_path_wires[7][2] ),
    .A2(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[7][3] ),
    .X(_08277_));
 sky130_fd_sc_hd__nand4_2 _15661_ (.A(\top_inst.grid_inst.data_path_wires[7][3] ),
    .B(_08139_),
    .C(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[3] ),
    .Y(_08278_));
 sky130_fd_sc_hd__a22o_1 _15662_ (.A1(_08163_),
    .A2(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[2] ),
    .B1(_08277_),
    .B2(_08278_),
    .X(_08279_));
 sky130_fd_sc_hd__nand4_2 _15663_ (.A(_08163_),
    .B(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[2] ),
    .C(_08277_),
    .D(_08278_),
    .Y(_08280_));
 sky130_fd_sc_hd__nand2_1 _15664_ (.A(_08279_),
    .B(_08280_),
    .Y(_08281_));
 sky130_fd_sc_hd__xnor2_1 _15665_ (.A(_08276_),
    .B(_08281_),
    .Y(_08282_));
 sky130_fd_sc_hd__xor2_1 _15666_ (.A(_08245_),
    .B(_08282_),
    .X(_08283_));
 sky130_fd_sc_hd__a21boi_1 _15667_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[5] ),
    .A2(_08250_),
    .B1_N(_08251_),
    .Y(_08284_));
 sky130_fd_sc_hd__a22o_1 _15668_ (.A1(\top_inst.grid_inst.data_path_wires[7][5] ),
    .A2(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[1] ),
    .B1(_08154_),
    .B2(\top_inst.grid_inst.data_path_wires[7][6] ),
    .X(_08285_));
 sky130_fd_sc_hd__nand4_1 _15669_ (.A(_08149_),
    .B(\top_inst.grid_inst.data_path_wires[7][5] ),
    .C(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[1] ),
    .D(_08154_),
    .Y(_08286_));
 sky130_fd_sc_hd__and3_1 _15670_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[6] ),
    .B(_08285_),
    .C(_08286_),
    .X(_08287_));
 sky130_fd_sc_hd__a21oi_1 _15671_ (.A1(_08285_),
    .A2(_08286_),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[6] ),
    .Y(_08288_));
 sky130_fd_sc_hd__a211o_1 _15672_ (.A1(_08241_),
    .A2(_08243_),
    .B1(_08287_),
    .C1(_08288_),
    .X(_08289_));
 sky130_fd_sc_hd__o211ai_1 _15673_ (.A1(_08287_),
    .A2(_08288_),
    .B1(_08241_),
    .C1(_08243_),
    .Y(_08290_));
 sky130_fd_sc_hd__and2_1 _15674_ (.A(_08289_),
    .B(_08290_),
    .X(_08291_));
 sky130_fd_sc_hd__xnor2_1 _15675_ (.A(_08284_),
    .B(_08291_),
    .Y(_08292_));
 sky130_fd_sc_hd__nand2_1 _15676_ (.A(_08283_),
    .B(_08292_),
    .Y(_08293_));
 sky130_fd_sc_hd__or2_1 _15677_ (.A(_08283_),
    .B(_08292_),
    .X(_08294_));
 sky130_fd_sc_hd__and2_1 _15678_ (.A(_08247_),
    .B(_08255_),
    .X(_08295_));
 sky130_fd_sc_hd__a21oi_1 _15679_ (.A1(_08293_),
    .A2(_08294_),
    .B1(_08295_),
    .Y(_08296_));
 sky130_fd_sc_hd__and3_1 _15680_ (.A(_08295_),
    .B(_08293_),
    .C(_08294_),
    .X(_08297_));
 sky130_fd_sc_hd__a211oi_2 _15681_ (.A1(_08272_),
    .A2(_08273_),
    .B1(_08296_),
    .C1(_08297_),
    .Y(_08298_));
 sky130_fd_sc_hd__o211a_1 _15682_ (.A1(_08296_),
    .A2(_08297_),
    .B1(_08272_),
    .C1(_08273_),
    .X(_08299_));
 sky130_fd_sc_hd__a211o_1 _15683_ (.A1(_08270_),
    .A2(_08271_),
    .B1(_08298_),
    .C1(_08299_),
    .X(_08300_));
 sky130_fd_sc_hd__o211ai_1 _15684_ (.A1(_08298_),
    .A2(_08299_),
    .B1(_08270_),
    .C1(_08271_),
    .Y(_08301_));
 sky130_fd_sc_hd__and3_1 _15685_ (.A(_08269_),
    .B(_08300_),
    .C(_08301_),
    .X(_08302_));
 sky130_fd_sc_hd__a21oi_1 _15686_ (.A1(_08300_),
    .A2(_08301_),
    .B1(_08269_),
    .Y(_08303_));
 sky130_fd_sc_hd__nor2_1 _15687_ (.A(_08302_),
    .B(_08303_),
    .Y(_08304_));
 sky130_fd_sc_hd__o31a_1 _15688_ (.A1(_08211_),
    .A2(_08233_),
    .A3(_08260_),
    .B1(_08264_),
    .X(_08305_));
 sky130_fd_sc_hd__xnor2_2 _15689_ (.A(_08304_),
    .B(_08305_),
    .Y(_08306_));
 sky130_fd_sc_hd__buf_8 _15690_ (.A(_05311_),
    .X(_08307_));
 sky130_fd_sc_hd__mux2_1 _15691_ (.A0(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[6] ),
    .A1(_08306_),
    .S(_08307_),
    .X(_08308_));
 sky130_fd_sc_hd__and2_1 _15692_ (.A(_08197_),
    .B(_08308_),
    .X(_08309_));
 sky130_fd_sc_hd__clkbuf_1 _15693_ (.A(_08309_),
    .X(_00505_));
 sky130_fd_sc_hd__nor2_1 _15694_ (.A(_08276_),
    .B(_08281_),
    .Y(_08310_));
 sky130_fd_sc_hd__nand2_1 _15695_ (.A(\top_inst.grid_inst.data_path_wires[7][1] ),
    .B(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[6] ),
    .Y(_08311_));
 sky130_fd_sc_hd__or2b_1 _15696_ (.A(\top_inst.grid_inst.data_path_wires[7][0] ),
    .B_N(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[7] ),
    .X(_08312_));
 sky130_fd_sc_hd__xnor2_1 _15697_ (.A(_08311_),
    .B(_08312_),
    .Y(_08313_));
 sky130_fd_sc_hd__nand2_1 _15698_ (.A(\top_inst.grid_inst.data_path_wires[7][2] ),
    .B(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[5] ),
    .Y(_08314_));
 sky130_fd_sc_hd__xnor2_1 _15699_ (.A(_08313_),
    .B(_08314_),
    .Y(_08315_));
 sky130_fd_sc_hd__xor2_1 _15700_ (.A(_08275_),
    .B(_08315_),
    .X(_08316_));
 sky130_fd_sc_hd__a22o_1 _15701_ (.A1(\top_inst.grid_inst.data_path_wires[7][3] ),
    .A2(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[7][4] ),
    .X(_08317_));
 sky130_fd_sc_hd__nand4_2 _15702_ (.A(\top_inst.grid_inst.data_path_wires[7][4] ),
    .B(\top_inst.grid_inst.data_path_wires[7][3] ),
    .C(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[3] ),
    .Y(_08318_));
 sky130_fd_sc_hd__a22o_1 _15703_ (.A1(_08147_),
    .A2(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[2] ),
    .B1(_08317_),
    .B2(_08318_),
    .X(_08319_));
 sky130_fd_sc_hd__nand4_2 _15704_ (.A(_08147_),
    .B(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[2] ),
    .C(_08317_),
    .D(_08318_),
    .Y(_08320_));
 sky130_fd_sc_hd__nand2_1 _15705_ (.A(_08319_),
    .B(_08320_),
    .Y(_08321_));
 sky130_fd_sc_hd__xnor2_1 _15706_ (.A(_08316_),
    .B(_08321_),
    .Y(_08322_));
 sky130_fd_sc_hd__xnor2_1 _15707_ (.A(_08310_),
    .B(_08322_),
    .Y(_08323_));
 sky130_fd_sc_hd__a21bo_1 _15708_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[6] ),
    .A2(_08285_),
    .B1_N(_08286_),
    .X(_08324_));
 sky130_fd_sc_hd__a22o_1 _15709_ (.A1(_08149_),
    .A2(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[1] ),
    .B1(_08154_),
    .B2(\top_inst.grid_inst.data_path_wires[7][7] ),
    .X(_08325_));
 sky130_fd_sc_hd__nand4_1 _15710_ (.A(\top_inst.grid_inst.data_path_wires[7][7] ),
    .B(_08149_),
    .C(_08157_),
    .D(_08154_),
    .Y(_08326_));
 sky130_fd_sc_hd__and3_1 _15711_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[7] ),
    .B(_08325_),
    .C(_08326_),
    .X(_08327_));
 sky130_fd_sc_hd__a21oi_1 _15712_ (.A1(_08325_),
    .A2(_08326_),
    .B1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[7] ),
    .Y(_08328_));
 sky130_fd_sc_hd__a211oi_1 _15713_ (.A1(_08278_),
    .A2(_08280_),
    .B1(_08327_),
    .C1(_08328_),
    .Y(_08329_));
 sky130_fd_sc_hd__o211a_1 _15714_ (.A1(_08327_),
    .A2(_08328_),
    .B1(_08278_),
    .C1(_08280_),
    .X(_08330_));
 sky130_fd_sc_hd__nor2_1 _15715_ (.A(_08329_),
    .B(_08330_),
    .Y(_08331_));
 sky130_fd_sc_hd__xnor2_2 _15716_ (.A(_08324_),
    .B(_08331_),
    .Y(_08332_));
 sky130_fd_sc_hd__xor2_1 _15717_ (.A(_08323_),
    .B(_08332_),
    .X(_08333_));
 sky130_fd_sc_hd__o21ai_1 _15718_ (.A1(_08245_),
    .A2(_08282_),
    .B1(_08293_),
    .Y(_08334_));
 sky130_fd_sc_hd__xnor2_1 _15719_ (.A(_08333_),
    .B(_08334_),
    .Y(_08335_));
 sky130_fd_sc_hd__or2b_1 _15720_ (.A(_08284_),
    .B_N(_08291_),
    .X(_08336_));
 sky130_fd_sc_hd__nand2_1 _15721_ (.A(_08289_),
    .B(_08336_),
    .Y(_08337_));
 sky130_fd_sc_hd__xnor2_1 _15722_ (.A(_08335_),
    .B(_08337_),
    .Y(_08338_));
 sky130_fd_sc_hd__nor2_1 _15723_ (.A(_08297_),
    .B(_08298_),
    .Y(_08339_));
 sky130_fd_sc_hd__xnor2_1 _15724_ (.A(_08338_),
    .B(_08339_),
    .Y(_08340_));
 sky130_fd_sc_hd__xnor2_1 _15725_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[7] ),
    .B(_08340_),
    .Y(_08341_));
 sky130_fd_sc_hd__xor2_1 _15726_ (.A(_08300_),
    .B(_08341_),
    .X(_08342_));
 sky130_fd_sc_hd__o21bai_2 _15727_ (.A1(_08303_),
    .A2(_08305_),
    .B1_N(_08302_),
    .Y(_08343_));
 sky130_fd_sc_hd__nor2_1 _15728_ (.A(_08342_),
    .B(_08343_),
    .Y(_08344_));
 sky130_fd_sc_hd__a21o_1 _15729_ (.A1(_08342_),
    .A2(_08343_),
    .B1(_06404_),
    .X(_08345_));
 sky130_fd_sc_hd__a2bb2o_1 _15730_ (.A1_N(_08344_),
    .A2_N(_08345_),
    .B1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[7] ),
    .B2(_07816_),
    .X(_08346_));
 sky130_fd_sc_hd__and2_1 _15731_ (.A(_08197_),
    .B(_08346_),
    .X(_08347_));
 sky130_fd_sc_hd__clkbuf_1 _15732_ (.A(_08347_),
    .X(_00506_));
 sky130_fd_sc_hd__nor2_1 _15733_ (.A(_08300_),
    .B(_08341_),
    .Y(_08348_));
 sky130_fd_sc_hd__a21o_1 _15734_ (.A1(_08342_),
    .A2(_08343_),
    .B1(_08348_),
    .X(_08349_));
 sky130_fd_sc_hd__or2b_1 _15735_ (.A(_08339_),
    .B_N(_08338_),
    .X(_08350_));
 sky130_fd_sc_hd__nand2_1 _15736_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[7] ),
    .B(_08340_),
    .Y(_08351_));
 sky130_fd_sc_hd__and4b_1 _15737_ (.A_N(\top_inst.grid_inst.data_path_wires[7][1] ),
    .B(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[7] ),
    .C(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[6] ),
    .D(\top_inst.grid_inst.data_path_wires[7][2] ),
    .X(_08352_));
 sky130_fd_sc_hd__inv_2 _15738_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[7] ),
    .Y(_08353_));
 sky130_fd_sc_hd__o2bb2a_1 _15739_ (.A1_N(\top_inst.grid_inst.data_path_wires[7][2] ),
    .A2_N(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[6] ),
    .B1(_08353_),
    .B2(\top_inst.grid_inst.data_path_wires[7][1] ),
    .X(_08354_));
 sky130_fd_sc_hd__nor2_2 _15740_ (.A(_08352_),
    .B(_08354_),
    .Y(_08355_));
 sky130_fd_sc_hd__nand2_2 _15741_ (.A(_08143_),
    .B(_08167_),
    .Y(_08356_));
 sky130_fd_sc_hd__xnor2_4 _15742_ (.A(_08355_),
    .B(_08356_),
    .Y(_08357_));
 sky130_fd_sc_hd__nor2_1 _15743_ (.A(_08313_),
    .B(_08314_),
    .Y(_08358_));
 sky130_fd_sc_hd__o21ba_1 _15744_ (.A1(_08311_),
    .A2(_08312_),
    .B1_N(_08358_),
    .X(_08359_));
 sky130_fd_sc_hd__xnor2_2 _15745_ (.A(_08357_),
    .B(_08359_),
    .Y(_08360_));
 sky130_fd_sc_hd__a22o_1 _15746_ (.A1(_08163_),
    .A2(_08164_),
    .B1(_08161_),
    .B2(_08147_),
    .X(_08361_));
 sky130_fd_sc_hd__nand4_4 _15747_ (.A(_08147_),
    .B(_08163_),
    .C(_08164_),
    .D(_08161_),
    .Y(_08362_));
 sky130_fd_sc_hd__a22o_1 _15748_ (.A1(_08149_),
    .A2(_08159_),
    .B1(_08361_),
    .B2(_08362_),
    .X(_08363_));
 sky130_fd_sc_hd__nand4_4 _15749_ (.A(_08150_),
    .B(_08159_),
    .C(_08361_),
    .D(_08362_),
    .Y(_08364_));
 sky130_fd_sc_hd__nand2_1 _15750_ (.A(_08363_),
    .B(_08364_),
    .Y(_08365_));
 sky130_fd_sc_hd__xnor2_1 _15751_ (.A(_08360_),
    .B(_08365_),
    .Y(_08366_));
 sky130_fd_sc_hd__and3_1 _15752_ (.A(_08316_),
    .B(_08319_),
    .C(_08320_),
    .X(_08367_));
 sky130_fd_sc_hd__o21ba_1 _15753_ (.A1(_08275_),
    .A2(_08315_),
    .B1_N(_08367_),
    .X(_08368_));
 sky130_fd_sc_hd__xnor2_1 _15754_ (.A(_08366_),
    .B(_08368_),
    .Y(_08369_));
 sky130_fd_sc_hd__and4_1 _15755_ (.A(_08152_),
    .B(_08150_),
    .C(_08157_),
    .D(_08155_),
    .X(_08370_));
 sky130_fd_sc_hd__o21ai_2 _15756_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[1] ),
    .A2(_08154_),
    .B1(\top_inst.grid_inst.data_path_wires[7][7] ),
    .Y(_08371_));
 sky130_fd_sc_hd__and3_1 _15757_ (.A(\top_inst.grid_inst.data_path_wires[7][7] ),
    .B(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[1] ),
    .C(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[0] ),
    .X(_08372_));
 sky130_fd_sc_hd__clkbuf_4 _15758_ (.A(_08372_),
    .X(_08373_));
 sky130_fd_sc_hd__nor2_4 _15759_ (.A(_08371_),
    .B(_08373_),
    .Y(_08374_));
 sky130_fd_sc_hd__xnor2_1 _15760_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[8] ),
    .B(_08374_),
    .Y(_08375_));
 sky130_fd_sc_hd__a21oi_1 _15761_ (.A1(_08318_),
    .A2(_08320_),
    .B1(_08375_),
    .Y(_08376_));
 sky130_fd_sc_hd__and3_1 _15762_ (.A(_08318_),
    .B(_08320_),
    .C(_08375_),
    .X(_08377_));
 sky130_fd_sc_hd__nor2_1 _15763_ (.A(_08376_),
    .B(_08377_),
    .Y(_08378_));
 sky130_fd_sc_hd__o21a_1 _15764_ (.A1(_08370_),
    .A2(_08327_),
    .B1(_08378_),
    .X(_08379_));
 sky130_fd_sc_hd__nor3_1 _15765_ (.A(_08370_),
    .B(_08327_),
    .C(_08378_),
    .Y(_08380_));
 sky130_fd_sc_hd__nor2_1 _15766_ (.A(_08379_),
    .B(_08380_),
    .Y(_08381_));
 sky130_fd_sc_hd__xnor2_1 _15767_ (.A(_08369_),
    .B(_08381_),
    .Y(_08382_));
 sky130_fd_sc_hd__nand2_1 _15768_ (.A(_08310_),
    .B(_08322_),
    .Y(_08383_));
 sky130_fd_sc_hd__o21a_1 _15769_ (.A1(_08323_),
    .A2(_08332_),
    .B1(_08383_),
    .X(_08384_));
 sky130_fd_sc_hd__xnor2_1 _15770_ (.A(_08382_),
    .B(_08384_),
    .Y(_08385_));
 sky130_fd_sc_hd__a21oi_2 _15771_ (.A1(_08324_),
    .A2(_08331_),
    .B1(_08329_),
    .Y(_08386_));
 sky130_fd_sc_hd__xnor2_1 _15772_ (.A(_08385_),
    .B(_08386_),
    .Y(_08387_));
 sky130_fd_sc_hd__and2b_1 _15773_ (.A_N(_08335_),
    .B(_08337_),
    .X(_08388_));
 sky130_fd_sc_hd__a21oi_1 _15774_ (.A1(_08333_),
    .A2(_08334_),
    .B1(_08388_),
    .Y(_08389_));
 sky130_fd_sc_hd__xnor2_1 _15775_ (.A(_08387_),
    .B(_08389_),
    .Y(_08390_));
 sky130_fd_sc_hd__a21o_1 _15776_ (.A1(_08350_),
    .A2(_08351_),
    .B1(_08390_),
    .X(_08391_));
 sky130_fd_sc_hd__nand3_1 _15777_ (.A(_08350_),
    .B(_08351_),
    .C(_08390_),
    .Y(_08392_));
 sky130_fd_sc_hd__and2_1 _15778_ (.A(_08391_),
    .B(_08392_),
    .X(_08393_));
 sky130_fd_sc_hd__xor2_1 _15779_ (.A(_08349_),
    .B(_08393_),
    .X(_08394_));
 sky130_fd_sc_hd__or2_1 _15780_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[8] ),
    .B(_07866_),
    .X(_08395_));
 sky130_fd_sc_hd__o211a_1 _15781_ (.A1(_06848_),
    .A2(_08394_),
    .B1(_08395_),
    .C1(_08166_),
    .X(_00507_));
 sky130_fd_sc_hd__nand2_1 _15782_ (.A(_08349_),
    .B(_08393_),
    .Y(_08396_));
 sky130_fd_sc_hd__or2_1 _15783_ (.A(_08387_),
    .B(_08389_),
    .X(_08397_));
 sky130_fd_sc_hd__and4b_1 _15784_ (.A_N(\top_inst.grid_inst.data_path_wires[7][2] ),
    .B(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[7] ),
    .C(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[6] ),
    .D(\top_inst.grid_inst.data_path_wires[7][3] ),
    .X(_08398_));
 sky130_fd_sc_hd__o2bb2a_1 _15785_ (.A1_N(\top_inst.grid_inst.data_path_wires[7][3] ),
    .A2_N(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[6] ),
    .B1(_08353_),
    .B2(\top_inst.grid_inst.data_path_wires[7][2] ),
    .X(_08399_));
 sky130_fd_sc_hd__nor2_1 _15786_ (.A(_08398_),
    .B(_08399_),
    .Y(_08400_));
 sky130_fd_sc_hd__nand2_1 _15787_ (.A(_08163_),
    .B(_08167_),
    .Y(_08401_));
 sky130_fd_sc_hd__xnor2_1 _15788_ (.A(_08400_),
    .B(_08401_),
    .Y(_08402_));
 sky130_fd_sc_hd__o21ba_1 _15789_ (.A1(_08354_),
    .A2(_08356_),
    .B1_N(_08352_),
    .X(_08403_));
 sky130_fd_sc_hd__xor2_1 _15790_ (.A(_08402_),
    .B(_08403_),
    .X(_08404_));
 sky130_fd_sc_hd__a22o_1 _15791_ (.A1(_08147_),
    .A2(_08164_),
    .B1(_08161_),
    .B2(_08149_),
    .X(_08405_));
 sky130_fd_sc_hd__and4_1 _15792_ (.A(\top_inst.grid_inst.data_path_wires[7][6] ),
    .B(\top_inst.grid_inst.data_path_wires[7][5] ),
    .C(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[3] ),
    .X(_08406_));
 sky130_fd_sc_hd__inv_2 _15793_ (.A(_08406_),
    .Y(_08407_));
 sky130_fd_sc_hd__and2_1 _15794_ (.A(_08405_),
    .B(_08407_),
    .X(_08408_));
 sky130_fd_sc_hd__nand2_4 _15795_ (.A(\top_inst.grid_inst.data_path_wires[7][7] ),
    .B(_08159_),
    .Y(_08409_));
 sky130_fd_sc_hd__xor2_1 _15796_ (.A(_08408_),
    .B(_08409_),
    .X(_08410_));
 sky130_fd_sc_hd__xor2_1 _15797_ (.A(_08404_),
    .B(_08410_),
    .X(_08411_));
 sky130_fd_sc_hd__inv_2 _15798_ (.A(_08359_),
    .Y(_08412_));
 sky130_fd_sc_hd__a32oi_4 _15799_ (.A1(_08360_),
    .A2(_08363_),
    .A3(_08364_),
    .B1(_08412_),
    .B2(_08357_),
    .Y(_08413_));
 sky130_fd_sc_hd__xnor2_1 _15800_ (.A(_08411_),
    .B(_08413_),
    .Y(_08414_));
 sky130_fd_sc_hd__a21o_1 _15801_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[8] ),
    .A2(_08374_),
    .B1(_08373_),
    .X(_08415_));
 sky130_fd_sc_hd__xnor2_1 _15802_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[9] ),
    .B(_08374_),
    .Y(_08416_));
 sky130_fd_sc_hd__a21oi_1 _15803_ (.A1(_08362_),
    .A2(_08364_),
    .B1(_08416_),
    .Y(_08417_));
 sky130_fd_sc_hd__and3_1 _15804_ (.A(_08362_),
    .B(_08364_),
    .C(_08416_),
    .X(_08418_));
 sky130_fd_sc_hd__nor2_1 _15805_ (.A(_08417_),
    .B(_08418_),
    .Y(_08419_));
 sky130_fd_sc_hd__xor2_1 _15806_ (.A(_08415_),
    .B(_08419_),
    .X(_08420_));
 sky130_fd_sc_hd__xnor2_1 _15807_ (.A(_08414_),
    .B(_08420_),
    .Y(_08421_));
 sky130_fd_sc_hd__and2b_1 _15808_ (.A_N(_08368_),
    .B(_08366_),
    .X(_08422_));
 sky130_fd_sc_hd__a21oi_1 _15809_ (.A1(_08369_),
    .A2(_08381_),
    .B1(_08422_),
    .Y(_08423_));
 sky130_fd_sc_hd__xnor2_1 _15810_ (.A(_08421_),
    .B(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__nor2_1 _15811_ (.A(_08376_),
    .B(_08379_),
    .Y(_08425_));
 sky130_fd_sc_hd__xnor2_1 _15812_ (.A(_08424_),
    .B(_08425_),
    .Y(_08426_));
 sky130_fd_sc_hd__or2_1 _15813_ (.A(_08382_),
    .B(_08384_),
    .X(_08427_));
 sky130_fd_sc_hd__o21a_1 _15814_ (.A1(_08385_),
    .A2(_08386_),
    .B1(_08427_),
    .X(_08428_));
 sky130_fd_sc_hd__nor2_1 _15815_ (.A(_08426_),
    .B(_08428_),
    .Y(_08429_));
 sky130_fd_sc_hd__and2_1 _15816_ (.A(_08426_),
    .B(_08428_),
    .X(_08430_));
 sky130_fd_sc_hd__or2_1 _15817_ (.A(_08429_),
    .B(_08430_),
    .X(_08431_));
 sky130_fd_sc_hd__xor2_2 _15818_ (.A(_08397_),
    .B(_08431_),
    .X(_08432_));
 sky130_fd_sc_hd__a21oi_1 _15819_ (.A1(_08391_),
    .A2(_08396_),
    .B1(_08432_),
    .Y(_08433_));
 sky130_fd_sc_hd__a31o_1 _15820_ (.A1(_08391_),
    .A2(_08396_),
    .A3(_08432_),
    .B1(_07439_),
    .X(_08434_));
 sky130_fd_sc_hd__o221a_1 _15821_ (.A1(net1086),
    .A2(_07048_),
    .B1(_08433_),
    .B2(_08434_),
    .C1(_07708_),
    .X(_00508_));
 sky130_fd_sc_hd__or2b_1 _15822_ (.A(_08403_),
    .B_N(_08402_),
    .X(_08435_));
 sky130_fd_sc_hd__o21a_1 _15823_ (.A1(_08404_),
    .A2(_08410_),
    .B1(_08435_),
    .X(_08436_));
 sky130_fd_sc_hd__and4b_1 _15824_ (.A_N(_08143_),
    .B(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[7] ),
    .C(_08169_),
    .D(_08163_),
    .X(_08437_));
 sky130_fd_sc_hd__o2bb2a_1 _15825_ (.A1_N(_08163_),
    .A2_N(_08169_),
    .B1(_08353_),
    .B2(_08143_),
    .X(_08438_));
 sky130_fd_sc_hd__nor2_1 _15826_ (.A(_08437_),
    .B(_08438_),
    .Y(_08439_));
 sky130_fd_sc_hd__nand2_1 _15827_ (.A(_08147_),
    .B(_08167_),
    .Y(_08440_));
 sky130_fd_sc_hd__xnor2_1 _15828_ (.A(_08439_),
    .B(_08440_),
    .Y(_08441_));
 sky130_fd_sc_hd__o21ba_1 _15829_ (.A1(_08399_),
    .A2(_08401_),
    .B1_N(_08398_),
    .X(_08442_));
 sky130_fd_sc_hd__xnor2_1 _15830_ (.A(_08441_),
    .B(_08442_),
    .Y(_08443_));
 sky130_fd_sc_hd__and3_1 _15831_ (.A(\top_inst.grid_inst.data_path_wires[7][7] ),
    .B(_08164_),
    .C(_08161_),
    .X(_08444_));
 sky130_fd_sc_hd__a22o_1 _15832_ (.A1(_08149_),
    .A2(_08164_),
    .B1(_08161_),
    .B2(\top_inst.grid_inst.data_path_wires[7][7] ),
    .X(_08445_));
 sky130_fd_sc_hd__a21bo_1 _15833_ (.A1(_08150_),
    .A2(_08444_),
    .B1_N(_08445_),
    .X(_08446_));
 sky130_fd_sc_hd__xor2_1 _15834_ (.A(_08409_),
    .B(_08446_),
    .X(_08447_));
 sky130_fd_sc_hd__xor2_1 _15835_ (.A(_08443_),
    .B(_08447_),
    .X(_08448_));
 sky130_fd_sc_hd__and2b_1 _15836_ (.A_N(_08436_),
    .B(_08448_),
    .X(_08449_));
 sky130_fd_sc_hd__and2b_1 _15837_ (.A_N(_08448_),
    .B(_08436_),
    .X(_08450_));
 sky130_fd_sc_hd__nor2_1 _15838_ (.A(_08449_),
    .B(_08450_),
    .Y(_08451_));
 sky130_fd_sc_hd__buf_4 _15839_ (.A(_08374_),
    .X(_08452_));
 sky130_fd_sc_hd__a21o_1 _15840_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[9] ),
    .A2(_08452_),
    .B1(_08373_),
    .X(_08453_));
 sky130_fd_sc_hd__a31o_1 _15841_ (.A1(_08152_),
    .A2(_08159_),
    .A3(_08405_),
    .B1(_08406_),
    .X(_08454_));
 sky130_fd_sc_hd__xnor2_1 _15842_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[10] ),
    .B(_08374_),
    .Y(_08455_));
 sky130_fd_sc_hd__xnor2_1 _15843_ (.A(_08454_),
    .B(_08455_),
    .Y(_08456_));
 sky130_fd_sc_hd__xor2_1 _15844_ (.A(_08453_),
    .B(_08456_),
    .X(_08457_));
 sky130_fd_sc_hd__xnor2_1 _15845_ (.A(_08451_),
    .B(_08457_),
    .Y(_08458_));
 sky130_fd_sc_hd__and2b_1 _15846_ (.A_N(_08413_),
    .B(_08411_),
    .X(_08459_));
 sky130_fd_sc_hd__a21oi_1 _15847_ (.A1(_08414_),
    .A2(_08420_),
    .B1(_08459_),
    .Y(_08460_));
 sky130_fd_sc_hd__xnor2_1 _15848_ (.A(_08458_),
    .B(_08460_),
    .Y(_08461_));
 sky130_fd_sc_hd__a21oi_1 _15849_ (.A1(_08415_),
    .A2(_08419_),
    .B1(_08417_),
    .Y(_08462_));
 sky130_fd_sc_hd__xnor2_1 _15850_ (.A(_08461_),
    .B(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__or2_1 _15851_ (.A(_08421_),
    .B(_08423_),
    .X(_08464_));
 sky130_fd_sc_hd__o21a_1 _15852_ (.A1(_08424_),
    .A2(_08425_),
    .B1(_08464_),
    .X(_08465_));
 sky130_fd_sc_hd__xor2_1 _15853_ (.A(_08463_),
    .B(_08465_),
    .X(_08466_));
 sky130_fd_sc_hd__and2_1 _15854_ (.A(_08429_),
    .B(_08466_),
    .X(_08467_));
 sky130_fd_sc_hd__nor2_1 _15855_ (.A(_08429_),
    .B(_08466_),
    .Y(_08468_));
 sky130_fd_sc_hd__nor2_1 _15856_ (.A(_08467_),
    .B(_08468_),
    .Y(_08469_));
 sky130_fd_sc_hd__a21oi_1 _15857_ (.A1(_08397_),
    .A2(_08391_),
    .B1(_08431_),
    .Y(_08470_));
 sky130_fd_sc_hd__a31o_1 _15858_ (.A1(_08349_),
    .A2(_08393_),
    .A3(_08432_),
    .B1(_08470_),
    .X(_08471_));
 sky130_fd_sc_hd__nand2_1 _15859_ (.A(_08469_),
    .B(_08471_),
    .Y(_08472_));
 sky130_fd_sc_hd__o21a_1 _15860_ (.A1(_08469_),
    .A2(_08471_),
    .B1(_08265_),
    .X(_08473_));
 sky130_fd_sc_hd__a22o_1 _15861_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[10] ),
    .A2(_08066_),
    .B1(_08472_),
    .B2(_08473_),
    .X(_08474_));
 sky130_fd_sc_hd__and2_1 _15862_ (.A(_08197_),
    .B(_08474_),
    .X(_08475_));
 sky130_fd_sc_hd__clkbuf_1 _15863_ (.A(_08475_),
    .X(_00509_));
 sky130_fd_sc_hd__inv_2 _15864_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[11] ),
    .Y(_08476_));
 sky130_fd_sc_hd__nor2_1 _15865_ (.A(_08463_),
    .B(_08465_),
    .Y(_08477_));
 sky130_fd_sc_hd__nor2_1 _15866_ (.A(_08458_),
    .B(_08460_),
    .Y(_08478_));
 sky130_fd_sc_hd__nor2_1 _15867_ (.A(_08461_),
    .B(_08462_),
    .Y(_08479_));
 sky130_fd_sc_hd__or2b_1 _15868_ (.A(_08442_),
    .B_N(_08441_),
    .X(_08480_));
 sky130_fd_sc_hd__nand2_1 _15869_ (.A(_08443_),
    .B(_08447_),
    .Y(_08481_));
 sky130_fd_sc_hd__o21ai_1 _15870_ (.A1(_08164_),
    .A2(_08161_),
    .B1(\top_inst.grid_inst.data_path_wires[7][7] ),
    .Y(_08482_));
 sky130_fd_sc_hd__nor2_2 _15871_ (.A(_08444_),
    .B(_08482_),
    .Y(_08483_));
 sky130_fd_sc_hd__xnor2_4 _15872_ (.A(_08409_),
    .B(_08483_),
    .Y(_08484_));
 sky130_fd_sc_hd__and4_1 _15873_ (.A(\top_inst.grid_inst.data_path_wires[7][5] ),
    .B(_08145_),
    .C(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[7] ),
    .D(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[6] ),
    .X(_08485_));
 sky130_fd_sc_hd__a22o_1 _15874_ (.A1(_08145_),
    .A2(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[7] ),
    .B1(_08169_),
    .B2(\top_inst.grid_inst.data_path_wires[7][5] ),
    .X(_08486_));
 sky130_fd_sc_hd__and2b_1 _15875_ (.A_N(_08485_),
    .B(_08486_),
    .X(_08487_));
 sky130_fd_sc_hd__nand2_1 _15876_ (.A(_08149_),
    .B(_08167_),
    .Y(_08488_));
 sky130_fd_sc_hd__xnor2_1 _15877_ (.A(_08487_),
    .B(_08488_),
    .Y(_08489_));
 sky130_fd_sc_hd__o21ba_1 _15878_ (.A1(_08438_),
    .A2(_08440_),
    .B1_N(_08437_),
    .X(_08490_));
 sky130_fd_sc_hd__xnor2_1 _15879_ (.A(_08489_),
    .B(_08490_),
    .Y(_08491_));
 sky130_fd_sc_hd__nand2_1 _15880_ (.A(_08484_),
    .B(_08491_),
    .Y(_08492_));
 sky130_fd_sc_hd__or2_1 _15881_ (.A(_08484_),
    .B(_08491_),
    .X(_08493_));
 sky130_fd_sc_hd__nand2_1 _15882_ (.A(_08492_),
    .B(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__a21oi_1 _15883_ (.A1(_08480_),
    .A2(_08481_),
    .B1(_08494_),
    .Y(_08495_));
 sky130_fd_sc_hd__nand3_1 _15884_ (.A(_08480_),
    .B(_08481_),
    .C(_08494_),
    .Y(_08496_));
 sky130_fd_sc_hd__or2b_1 _15885_ (.A(_08495_),
    .B_N(_08496_),
    .X(_08497_));
 sky130_fd_sc_hd__a21o_1 _15886_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[10] ),
    .A2(_08452_),
    .B1(_08373_),
    .X(_08498_));
 sky130_fd_sc_hd__a32o_1 _15887_ (.A1(_08152_),
    .A2(_08159_),
    .A3(_08445_),
    .B1(_08444_),
    .B2(_08150_),
    .X(_08499_));
 sky130_fd_sc_hd__xnor2_1 _15888_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[11] ),
    .B(_08374_),
    .Y(_08500_));
 sky130_fd_sc_hd__xnor2_1 _15889_ (.A(_08499_),
    .B(_08500_),
    .Y(_08501_));
 sky130_fd_sc_hd__xor2_1 _15890_ (.A(_08498_),
    .B(_08501_),
    .X(_08502_));
 sky130_fd_sc_hd__xnor2_1 _15891_ (.A(_08497_),
    .B(_08502_),
    .Y(_08503_));
 sky130_fd_sc_hd__a21o_1 _15892_ (.A1(_08451_),
    .A2(_08457_),
    .B1(_08449_),
    .X(_08504_));
 sky130_fd_sc_hd__xnor2_1 _15893_ (.A(_08503_),
    .B(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__or2b_1 _15894_ (.A(_08455_),
    .B_N(_08454_),
    .X(_08506_));
 sky130_fd_sc_hd__a21bo_1 _15895_ (.A1(_08453_),
    .A2(_08456_),
    .B1_N(_08506_),
    .X(_08507_));
 sky130_fd_sc_hd__xnor2_1 _15896_ (.A(_08505_),
    .B(_08507_),
    .Y(_08508_));
 sky130_fd_sc_hd__o21ai_2 _15897_ (.A1(_08478_),
    .A2(_08479_),
    .B1(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__or3_1 _15898_ (.A(_08478_),
    .B(_08479_),
    .C(_08508_),
    .X(_08510_));
 sky130_fd_sc_hd__and2_1 _15899_ (.A(_08509_),
    .B(_08510_),
    .X(_08511_));
 sky130_fd_sc_hd__xnor2_1 _15900_ (.A(_08477_),
    .B(_08511_),
    .Y(_08512_));
 sky130_fd_sc_hd__a21oi_1 _15901_ (.A1(_08469_),
    .A2(_08471_),
    .B1(_08467_),
    .Y(_08513_));
 sky130_fd_sc_hd__xnor2_1 _15902_ (.A(_08512_),
    .B(_08513_),
    .Y(_08514_));
 sky130_fd_sc_hd__mux2_1 _15903_ (.A0(_08476_),
    .A1(_08514_),
    .S(_05335_),
    .X(_08515_));
 sky130_fd_sc_hd__nor2_1 _15904_ (.A(_05632_),
    .B(_08515_),
    .Y(_00510_));
 sky130_fd_sc_hd__or2b_1 _15905_ (.A(_08490_),
    .B_N(_08489_),
    .X(_08516_));
 sky130_fd_sc_hd__nand2_2 _15906_ (.A(_08152_),
    .B(_08167_),
    .Y(_08517_));
 sky130_fd_sc_hd__nor2_1 _15907_ (.A(_08147_),
    .B(_08353_),
    .Y(_08518_));
 sky130_fd_sc_hd__and3_1 _15908_ (.A(_08149_),
    .B(_08169_),
    .C(_08518_),
    .X(_08519_));
 sky130_fd_sc_hd__a21oi_1 _15909_ (.A1(_08149_),
    .A2(_08169_),
    .B1(_08518_),
    .Y(_08520_));
 sky130_fd_sc_hd__or2_1 _15910_ (.A(_08519_),
    .B(_08520_),
    .X(_08521_));
 sky130_fd_sc_hd__xor2_1 _15911_ (.A(_08517_),
    .B(_08521_),
    .X(_08522_));
 sky130_fd_sc_hd__a31o_1 _15912_ (.A1(_08150_),
    .A2(_08167_),
    .A3(_08486_),
    .B1(_08485_),
    .X(_08523_));
 sky130_fd_sc_hd__xor2_1 _15913_ (.A(_08522_),
    .B(_08523_),
    .X(_08524_));
 sky130_fd_sc_hd__nand2_1 _15914_ (.A(_08484_),
    .B(_08524_),
    .Y(_08525_));
 sky130_fd_sc_hd__or2_1 _15915_ (.A(_08484_),
    .B(_08524_),
    .X(_08526_));
 sky130_fd_sc_hd__nand2_1 _15916_ (.A(_08525_),
    .B(_08526_),
    .Y(_08527_));
 sky130_fd_sc_hd__a21o_1 _15917_ (.A1(_08516_),
    .A2(_08492_),
    .B1(_08527_),
    .X(_08528_));
 sky130_fd_sc_hd__nand3_1 _15918_ (.A(_08516_),
    .B(_08492_),
    .C(_08527_),
    .Y(_08529_));
 sky130_fd_sc_hd__nand2_2 _15919_ (.A(_08528_),
    .B(_08529_),
    .Y(_08530_));
 sky130_fd_sc_hd__a21o_1 _15920_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[11] ),
    .A2(_08452_),
    .B1(_08373_),
    .X(_08531_));
 sky130_fd_sc_hd__o21ba_2 _15921_ (.A1(_08409_),
    .A2(_08482_),
    .B1_N(_08444_),
    .X(_08532_));
 sky130_fd_sc_hd__xnor2_1 _15922_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[12] ),
    .B(_08374_),
    .Y(_08533_));
 sky130_fd_sc_hd__nor2_1 _15923_ (.A(_08532_),
    .B(_08533_),
    .Y(_08534_));
 sky130_fd_sc_hd__and2_1 _15924_ (.A(_08532_),
    .B(_08533_),
    .X(_08535_));
 sky130_fd_sc_hd__nor2_1 _15925_ (.A(_08534_),
    .B(_08535_),
    .Y(_08536_));
 sky130_fd_sc_hd__xnor2_2 _15926_ (.A(_08531_),
    .B(_08536_),
    .Y(_08537_));
 sky130_fd_sc_hd__xor2_2 _15927_ (.A(_08530_),
    .B(_08537_),
    .X(_08538_));
 sky130_fd_sc_hd__a21o_1 _15928_ (.A1(_08496_),
    .A2(_08502_),
    .B1(_08495_),
    .X(_08539_));
 sky130_fd_sc_hd__xnor2_2 _15929_ (.A(_08538_),
    .B(_08539_),
    .Y(_08540_));
 sky130_fd_sc_hd__or2b_1 _15930_ (.A(_08500_),
    .B_N(_08499_),
    .X(_08541_));
 sky130_fd_sc_hd__a21bo_1 _15931_ (.A1(_08498_),
    .A2(_08501_),
    .B1_N(_08541_),
    .X(_08542_));
 sky130_fd_sc_hd__xnor2_2 _15932_ (.A(_08540_),
    .B(_08542_),
    .Y(_08543_));
 sky130_fd_sc_hd__or2b_1 _15933_ (.A(_08505_),
    .B_N(_08507_),
    .X(_08544_));
 sky130_fd_sc_hd__a21bo_1 _15934_ (.A1(_08503_),
    .A2(_08504_),
    .B1_N(_08544_),
    .X(_08545_));
 sky130_fd_sc_hd__and2_1 _15935_ (.A(_08543_),
    .B(_08545_),
    .X(_08546_));
 sky130_fd_sc_hd__nor2_1 _15936_ (.A(_08543_),
    .B(_08545_),
    .Y(_08547_));
 sky130_fd_sc_hd__nor2_1 _15937_ (.A(_08546_),
    .B(_08547_),
    .Y(_08548_));
 sky130_fd_sc_hd__xor2_2 _15938_ (.A(_08509_),
    .B(_08548_),
    .X(_08549_));
 sky130_fd_sc_hd__nand2_1 _15939_ (.A(_08477_),
    .B(_08511_),
    .Y(_08550_));
 sky130_fd_sc_hd__o21a_1 _15940_ (.A1(_08512_),
    .A2(_08513_),
    .B1(_08550_),
    .X(_08551_));
 sky130_fd_sc_hd__nor2_1 _15941_ (.A(_08549_),
    .B(_08551_),
    .Y(_08552_));
 sky130_fd_sc_hd__a21o_1 _15942_ (.A1(_08549_),
    .A2(_08551_),
    .B1(_06404_),
    .X(_08553_));
 sky130_fd_sc_hd__a2bb2o_1 _15943_ (.A1_N(_08552_),
    .A2_N(_08553_),
    .B1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[12] ),
    .B2(_07816_),
    .X(_08554_));
 sky130_fd_sc_hd__and2_1 _15944_ (.A(_08197_),
    .B(_08554_),
    .X(_08555_));
 sky130_fd_sc_hd__clkbuf_1 _15945_ (.A(_08555_),
    .X(_00511_));
 sky130_fd_sc_hd__nand2_1 _15946_ (.A(net1054),
    .B(_05403_),
    .Y(_08556_));
 sky130_fd_sc_hd__nand2_1 _15947_ (.A(_08522_),
    .B(_08523_),
    .Y(_08557_));
 sky130_fd_sc_hd__nand2_1 _15948_ (.A(_08152_),
    .B(_08169_),
    .Y(_08558_));
 sky130_fd_sc_hd__o21a_1 _15949_ (.A1(_08150_),
    .A2(_08353_),
    .B1(_08558_),
    .X(_08559_));
 sky130_fd_sc_hd__nor3_1 _15950_ (.A(_08150_),
    .B(_08353_),
    .C(_08558_),
    .Y(_08560_));
 sky130_fd_sc_hd__nor2_1 _15951_ (.A(_08559_),
    .B(_08560_),
    .Y(_08561_));
 sky130_fd_sc_hd__xnor2_1 _15952_ (.A(_08517_),
    .B(_08561_),
    .Y(_08562_));
 sky130_fd_sc_hd__o21ba_1 _15953_ (.A1(_08517_),
    .A2(_08520_),
    .B1_N(_08519_),
    .X(_08563_));
 sky130_fd_sc_hd__xnor2_1 _15954_ (.A(_08562_),
    .B(_08563_),
    .Y(_08564_));
 sky130_fd_sc_hd__nand2_1 _15955_ (.A(_08484_),
    .B(_08564_),
    .Y(_08565_));
 sky130_fd_sc_hd__or2_1 _15956_ (.A(_08484_),
    .B(_08564_),
    .X(_08566_));
 sky130_fd_sc_hd__nand2_1 _15957_ (.A(_08565_),
    .B(_08566_),
    .Y(_08567_));
 sky130_fd_sc_hd__a21o_1 _15958_ (.A1(_08557_),
    .A2(_08525_),
    .B1(_08567_),
    .X(_08568_));
 sky130_fd_sc_hd__nand3_1 _15959_ (.A(_08557_),
    .B(_08525_),
    .C(_08567_),
    .Y(_08569_));
 sky130_fd_sc_hd__a21o_1 _15960_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[12] ),
    .A2(_08452_),
    .B1(_08373_),
    .X(_08570_));
 sky130_fd_sc_hd__xnor2_1 _15961_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[13] ),
    .B(_08452_),
    .Y(_08571_));
 sky130_fd_sc_hd__nor2_1 _15962_ (.A(_08532_),
    .B(_08571_),
    .Y(_08572_));
 sky130_fd_sc_hd__and2_1 _15963_ (.A(_08532_),
    .B(_08571_),
    .X(_08573_));
 sky130_fd_sc_hd__nor2_1 _15964_ (.A(_08572_),
    .B(_08573_),
    .Y(_08574_));
 sky130_fd_sc_hd__xor2_1 _15965_ (.A(_08570_),
    .B(_08574_),
    .X(_08575_));
 sky130_fd_sc_hd__and3_1 _15966_ (.A(_08568_),
    .B(_08569_),
    .C(_08575_),
    .X(_08576_));
 sky130_fd_sc_hd__a21oi_1 _15967_ (.A1(_08568_),
    .A2(_08569_),
    .B1(_08575_),
    .Y(_08577_));
 sky130_fd_sc_hd__nor2_1 _15968_ (.A(_08576_),
    .B(_08577_),
    .Y(_08578_));
 sky130_fd_sc_hd__o21ai_2 _15969_ (.A1(_08530_),
    .A2(_08537_),
    .B1(_08528_),
    .Y(_08579_));
 sky130_fd_sc_hd__xnor2_1 _15970_ (.A(_08578_),
    .B(_08579_),
    .Y(_08580_));
 sky130_fd_sc_hd__a21o_1 _15971_ (.A1(_08531_),
    .A2(_08536_),
    .B1(_08534_),
    .X(_08581_));
 sky130_fd_sc_hd__xnor2_1 _15972_ (.A(_08580_),
    .B(_08581_),
    .Y(_08582_));
 sky130_fd_sc_hd__or2b_1 _15973_ (.A(_08540_),
    .B_N(_08542_),
    .X(_08583_));
 sky130_fd_sc_hd__a21bo_1 _15974_ (.A1(_08538_),
    .A2(_08539_),
    .B1_N(_08583_),
    .X(_08584_));
 sky130_fd_sc_hd__nand2_1 _15975_ (.A(_08582_),
    .B(_08584_),
    .Y(_08585_));
 sky130_fd_sc_hd__or2_1 _15976_ (.A(_08582_),
    .B(_08584_),
    .X(_08586_));
 sky130_fd_sc_hd__and2_1 _15977_ (.A(_08585_),
    .B(_08586_),
    .X(_08587_));
 sky130_fd_sc_hd__xor2_1 _15978_ (.A(_08546_),
    .B(_08587_),
    .X(_08588_));
 sky130_fd_sc_hd__and2b_1 _15979_ (.A_N(_08509_),
    .B(_08548_),
    .X(_08589_));
 sky130_fd_sc_hd__o21bai_2 _15980_ (.A1(_08549_),
    .A2(_08551_),
    .B1_N(_08589_),
    .Y(_08590_));
 sky130_fd_sc_hd__a21oi_1 _15981_ (.A1(_08588_),
    .A2(_08590_),
    .B1(_06734_),
    .Y(_08591_));
 sky130_fd_sc_hd__o21ai_1 _15982_ (.A1(_08588_),
    .A2(_08590_),
    .B1(_08591_),
    .Y(_08592_));
 sky130_fd_sc_hd__a21oi_1 _15983_ (.A1(_08556_),
    .A2(_08592_),
    .B1(_05440_),
    .Y(_00512_));
 sky130_fd_sc_hd__a21oi_1 _15984_ (.A1(_08557_),
    .A2(_08525_),
    .B1(_08567_),
    .Y(_08593_));
 sky130_fd_sc_hd__or2b_1 _15985_ (.A(_08563_),
    .B_N(_08562_),
    .X(_08594_));
 sky130_fd_sc_hd__and3_1 _15986_ (.A(_08152_),
    .B(_08169_),
    .C(_08167_),
    .X(_08595_));
 sky130_fd_sc_hd__o21ba_1 _15987_ (.A1(_08517_),
    .A2(_08559_),
    .B1_N(_08560_),
    .X(_08596_));
 sky130_fd_sc_hd__o21a_1 _15988_ (.A1(_08152_),
    .A2(_08353_),
    .B1(_08558_),
    .X(_08597_));
 sky130_fd_sc_hd__a2bb2o_1 _15989_ (.A1_N(_08595_),
    .A2_N(_08596_),
    .B1(_08517_),
    .B2(_08597_),
    .X(_08598_));
 sky130_fd_sc_hd__xor2_1 _15990_ (.A(_08484_),
    .B(_08598_),
    .X(_08599_));
 sky130_fd_sc_hd__a21oi_1 _15991_ (.A1(_08594_),
    .A2(_08565_),
    .B1(_08599_),
    .Y(_08600_));
 sky130_fd_sc_hd__nand3_1 _15992_ (.A(_08594_),
    .B(_08565_),
    .C(_08599_),
    .Y(_08601_));
 sky130_fd_sc_hd__or2b_1 _15993_ (.A(_08600_),
    .B_N(_08601_),
    .X(_08602_));
 sky130_fd_sc_hd__a21oi_1 _15994_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[13] ),
    .A2(_08452_),
    .B1(_08373_),
    .Y(_08603_));
 sky130_fd_sc_hd__xnor2_1 _15995_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[14] ),
    .B(_08452_),
    .Y(_08604_));
 sky130_fd_sc_hd__nor2_1 _15996_ (.A(_08532_),
    .B(_08604_),
    .Y(_08605_));
 sky130_fd_sc_hd__and2_1 _15997_ (.A(_08532_),
    .B(_08604_),
    .X(_08606_));
 sky130_fd_sc_hd__nor2_1 _15998_ (.A(_08605_),
    .B(_08606_),
    .Y(_08607_));
 sky130_fd_sc_hd__xnor2_1 _15999_ (.A(_08603_),
    .B(_08607_),
    .Y(_08608_));
 sky130_fd_sc_hd__xnor2_1 _16000_ (.A(_08602_),
    .B(_08608_),
    .Y(_08609_));
 sky130_fd_sc_hd__o21ai_1 _16001_ (.A1(_08593_),
    .A2(_08576_),
    .B1(_08609_),
    .Y(_08610_));
 sky130_fd_sc_hd__or3_1 _16002_ (.A(_08593_),
    .B(_08576_),
    .C(_08609_),
    .X(_08611_));
 sky130_fd_sc_hd__nand2_1 _16003_ (.A(_08610_),
    .B(_08611_),
    .Y(_08612_));
 sky130_fd_sc_hd__a21oi_2 _16004_ (.A1(_08570_),
    .A2(_08574_),
    .B1(_08572_),
    .Y(_08613_));
 sky130_fd_sc_hd__xnor2_2 _16005_ (.A(_08612_),
    .B(_08613_),
    .Y(_08614_));
 sky130_fd_sc_hd__or2b_1 _16006_ (.A(_08580_),
    .B_N(_08581_),
    .X(_08615_));
 sky130_fd_sc_hd__a21boi_2 _16007_ (.A1(_08578_),
    .A2(_08579_),
    .B1_N(_08615_),
    .Y(_08616_));
 sky130_fd_sc_hd__xnor2_1 _16008_ (.A(_08614_),
    .B(_08616_),
    .Y(_08617_));
 sky130_fd_sc_hd__nor2_1 _16009_ (.A(_08585_),
    .B(_08617_),
    .Y(_08618_));
 sky130_fd_sc_hd__and2_1 _16010_ (.A(_08585_),
    .B(_08617_),
    .X(_08619_));
 sky130_fd_sc_hd__nor2_2 _16011_ (.A(_08618_),
    .B(_08619_),
    .Y(_08620_));
 sky130_fd_sc_hd__a32o_2 _16012_ (.A1(_08543_),
    .A2(_08545_),
    .A3(_08587_),
    .B1(_08588_),
    .B2(_08590_),
    .X(_08621_));
 sky130_fd_sc_hd__nand2_1 _16013_ (.A(_08620_),
    .B(_08621_),
    .Y(_08622_));
 sky130_fd_sc_hd__o21a_1 _16014_ (.A1(_08620_),
    .A2(_08621_),
    .B1(_08265_),
    .X(_08623_));
 sky130_fd_sc_hd__a22o_1 _16015_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[14] ),
    .A2(_08066_),
    .B1(_08622_),
    .B2(_08623_),
    .X(_08624_));
 sky130_fd_sc_hd__and2_1 _16016_ (.A(_08197_),
    .B(_08624_),
    .X(_08625_));
 sky130_fd_sc_hd__clkbuf_1 _16017_ (.A(_08625_),
    .X(_00513_));
 sky130_fd_sc_hd__and2_1 _16018_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[15] ),
    .B(_07576_),
    .X(_08626_));
 sky130_fd_sc_hd__a21oi_1 _16019_ (.A1(_08601_),
    .A2(_08608_),
    .B1(_08600_),
    .Y(_08627_));
 sky130_fd_sc_hd__and2b_1 _16020_ (.A_N(_08484_),
    .B(_08598_),
    .X(_08628_));
 sky130_fd_sc_hd__a21o_1 _16021_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[14] ),
    .A2(_08452_),
    .B1(_08373_),
    .X(_08629_));
 sky130_fd_sc_hd__xnor2_2 _16022_ (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[15] ),
    .B(_08452_),
    .Y(_08630_));
 sky130_fd_sc_hd__xnor2_1 _16023_ (.A(_08532_),
    .B(_08630_),
    .Y(_08631_));
 sky130_fd_sc_hd__xnor2_1 _16024_ (.A(_08629_),
    .B(_08631_),
    .Y(_08632_));
 sky130_fd_sc_hd__or2_1 _16025_ (.A(_08628_),
    .B(_08632_),
    .X(_08633_));
 sky130_fd_sc_hd__nand2_1 _16026_ (.A(_08628_),
    .B(_08632_),
    .Y(_08634_));
 sky130_fd_sc_hd__and2_1 _16027_ (.A(_08633_),
    .B(_08634_),
    .X(_08635_));
 sky130_fd_sc_hd__xnor2_1 _16028_ (.A(_08627_),
    .B(_08635_),
    .Y(_08636_));
 sky130_fd_sc_hd__o21ba_1 _16029_ (.A1(_08603_),
    .A2(_08606_),
    .B1_N(_08605_),
    .X(_08637_));
 sky130_fd_sc_hd__xnor2_1 _16030_ (.A(_08636_),
    .B(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__o21a_1 _16031_ (.A1(_08612_),
    .A2(_08613_),
    .B1(_08610_),
    .X(_08639_));
 sky130_fd_sc_hd__or2_1 _16032_ (.A(_08638_),
    .B(_08639_),
    .X(_08640_));
 sky130_fd_sc_hd__nand2_1 _16033_ (.A(_08638_),
    .B(_08639_),
    .Y(_08641_));
 sky130_fd_sc_hd__and4bb_1 _16034_ (.A_N(_08614_),
    .B_N(_08616_),
    .C(_08640_),
    .D(_08641_),
    .X(_08642_));
 sky130_fd_sc_hd__and2_1 _16035_ (.A(_08640_),
    .B(_08641_),
    .X(_08643_));
 sky130_fd_sc_hd__o21ba_1 _16036_ (.A1(_08614_),
    .A2(_08616_),
    .B1_N(_08643_),
    .X(_08644_));
 sky130_fd_sc_hd__a21oi_1 _16037_ (.A1(_08620_),
    .A2(_08621_),
    .B1(_08618_),
    .Y(_08645_));
 sky130_fd_sc_hd__nor2_1 _16038_ (.A(_08642_),
    .B(_08644_),
    .Y(_08646_));
 sky130_fd_sc_hd__a211o_1 _16039_ (.A1(_08620_),
    .A2(_08621_),
    .B1(_08646_),
    .C1(_08618_),
    .X(_08647_));
 sky130_fd_sc_hd__o311a_1 _16040_ (.A1(_08642_),
    .A2(_08644_),
    .A3(_08645_),
    .B1(_08647_),
    .C1(_05313_),
    .X(_08648_));
 sky130_fd_sc_hd__o21a_1 _16041_ (.A1(_08626_),
    .A2(_08648_),
    .B1(_04870_),
    .X(_00514_));
 sky130_fd_sc_hd__or2_1 _16042_ (.A(_08627_),
    .B(_08635_),
    .X(_08649_));
 sky130_fd_sc_hd__o21a_1 _16043_ (.A1(_08636_),
    .A2(_08637_),
    .B1(_08649_),
    .X(_08650_));
 sky130_fd_sc_hd__xnor2_1 _16044_ (.A(_08633_),
    .B(_08650_),
    .Y(_08651_));
 sky130_fd_sc_hd__a21o_1 _16045_ (.A1(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[15] ),
    .A2(_08452_),
    .B1(_08373_),
    .X(_08652_));
 sky130_fd_sc_hd__o21a_1 _16046_ (.A1(_08532_),
    .A2(_08630_),
    .B1(_08629_),
    .X(_08653_));
 sky130_fd_sc_hd__a21oi_1 _16047_ (.A1(_08532_),
    .A2(_08630_),
    .B1(_08653_),
    .Y(_08654_));
 sky130_fd_sc_hd__xnor2_1 _16048_ (.A(_08640_),
    .B(_08654_),
    .Y(_08655_));
 sky130_fd_sc_hd__xnor2_1 _16049_ (.A(_08652_),
    .B(_08655_),
    .Y(_08656_));
 sky130_fd_sc_hd__xnor2_1 _16050_ (.A(_08651_),
    .B(_08656_),
    .Y(_08657_));
 sky130_fd_sc_hd__nor2_1 _16051_ (.A(_08642_),
    .B(_08657_),
    .Y(_08658_));
 sky130_fd_sc_hd__o31a_1 _16052_ (.A1(_08642_),
    .A2(_08644_),
    .A3(_08645_),
    .B1(_08658_),
    .X(_08659_));
 sky130_fd_sc_hd__or2_1 _16053_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[16] ),
    .B(_07866_),
    .X(_08660_));
 sky130_fd_sc_hd__o211a_1 _16054_ (.A1(_06848_),
    .A2(_08659_),
    .B1(_08660_),
    .C1(_08166_),
    .X(_00515_));
 sky130_fd_sc_hd__buf_2 _16055_ (.A(\top_inst.grid_inst.data_path_wires[8][0] ),
    .X(_08661_));
 sky130_fd_sc_hd__or2_1 _16056_ (.A(_08661_),
    .B(_08140_),
    .X(_08662_));
 sky130_fd_sc_hd__o211a_1 _16057_ (.A1(_08135_),
    .A2(_06634_),
    .B1(_08662_),
    .C1(_08166_),
    .X(_00516_));
 sky130_fd_sc_hd__buf_4 _16058_ (.A(_05177_),
    .X(_08663_));
 sky130_fd_sc_hd__buf_2 _16059_ (.A(\top_inst.grid_inst.data_path_wires[8][1] ),
    .X(_08664_));
 sky130_fd_sc_hd__or2_1 _16060_ (.A(_08664_),
    .B(_08140_),
    .X(_08665_));
 sky130_fd_sc_hd__buf_2 _16061_ (.A(_07617_),
    .X(_08666_));
 sky130_fd_sc_hd__o211a_1 _16062_ (.A1(_08137_),
    .A2(_08663_),
    .B1(_08665_),
    .C1(_08666_),
    .X(_00517_));
 sky130_fd_sc_hd__clkbuf_4 _16063_ (.A(\top_inst.grid_inst.data_path_wires[8][2] ),
    .X(_08667_));
 sky130_fd_sc_hd__or2_1 _16064_ (.A(_08667_),
    .B(_08140_),
    .X(_08668_));
 sky130_fd_sc_hd__o211a_1 _16065_ (.A1(_08139_),
    .A2(_08663_),
    .B1(_08668_),
    .C1(_08666_),
    .X(_00518_));
 sky130_fd_sc_hd__clkbuf_4 _16066_ (.A(\top_inst.grid_inst.data_path_wires[8][3] ),
    .X(_08669_));
 sky130_fd_sc_hd__or2_1 _16067_ (.A(_08669_),
    .B(_08140_),
    .X(_08670_));
 sky130_fd_sc_hd__o211a_1 _16068_ (.A1(_08143_),
    .A2(_08663_),
    .B1(_08670_),
    .C1(_08666_),
    .X(_00519_));
 sky130_fd_sc_hd__clkbuf_4 _16069_ (.A(\top_inst.grid_inst.data_path_wires[8][4] ),
    .X(_08671_));
 sky130_fd_sc_hd__or2_1 _16070_ (.A(_08671_),
    .B(_08140_),
    .X(_08672_));
 sky130_fd_sc_hd__o211a_1 _16071_ (.A1(_08163_),
    .A2(_08663_),
    .B1(_08672_),
    .C1(_08666_),
    .X(_00520_));
 sky130_fd_sc_hd__clkbuf_4 _16072_ (.A(\top_inst.grid_inst.data_path_wires[8][5] ),
    .X(_08673_));
 sky130_fd_sc_hd__clkbuf_4 _16073_ (.A(_06619_),
    .X(_08674_));
 sky130_fd_sc_hd__or2_1 _16074_ (.A(_08673_),
    .B(_08674_),
    .X(_08675_));
 sky130_fd_sc_hd__o211a_1 _16075_ (.A1(_08147_),
    .A2(_08663_),
    .B1(_08675_),
    .C1(_08666_),
    .X(_00521_));
 sky130_fd_sc_hd__buf_2 _16076_ (.A(\top_inst.grid_inst.data_path_wires[8][6] ),
    .X(_08676_));
 sky130_fd_sc_hd__clkbuf_4 _16077_ (.A(_08676_),
    .X(_08677_));
 sky130_fd_sc_hd__or2_1 _16078_ (.A(_08677_),
    .B(_08674_),
    .X(_08678_));
 sky130_fd_sc_hd__o211a_1 _16079_ (.A1(_08150_),
    .A2(_08663_),
    .B1(_08678_),
    .C1(_08666_),
    .X(_00522_));
 sky130_fd_sc_hd__clkbuf_4 _16080_ (.A(\top_inst.grid_inst.data_path_wires[8][7] ),
    .X(_08679_));
 sky130_fd_sc_hd__or2_1 _16081_ (.A(_08679_),
    .B(_08674_),
    .X(_08680_));
 sky130_fd_sc_hd__o211a_1 _16082_ (.A1(_08152_),
    .A2(_08663_),
    .B1(_08680_),
    .C1(_08666_),
    .X(_00523_));
 sky130_fd_sc_hd__clkbuf_4 _16083_ (.A(_05755_),
    .X(_08681_));
 sky130_fd_sc_hd__buf_2 _16084_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[0] ),
    .X(_08682_));
 sky130_fd_sc_hd__buf_2 _16085_ (.A(_08682_),
    .X(_08683_));
 sky130_fd_sc_hd__buf_2 _16086_ (.A(_05772_),
    .X(_08684_));
 sky130_fd_sc_hd__or2_1 _16087_ (.A(_08683_),
    .B(_08684_),
    .X(_08685_));
 sky130_fd_sc_hd__o211a_1 _16088_ (.A1(_08661_),
    .A2(_08681_),
    .B1(_08685_),
    .C1(_08666_),
    .X(_00524_));
 sky130_fd_sc_hd__buf_2 _16089_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[1] ),
    .X(_08686_));
 sky130_fd_sc_hd__or2_1 _16090_ (.A(_08686_),
    .B(_08684_),
    .X(_08687_));
 sky130_fd_sc_hd__o211a_1 _16091_ (.A1(_08664_),
    .A2(_08681_),
    .B1(_08687_),
    .C1(_08666_),
    .X(_00525_));
 sky130_fd_sc_hd__buf_4 _16092_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[2] ),
    .X(_08688_));
 sky130_fd_sc_hd__or2_1 _16093_ (.A(_08688_),
    .B(_08684_),
    .X(_08689_));
 sky130_fd_sc_hd__o211a_1 _16094_ (.A1(_08667_),
    .A2(_08681_),
    .B1(_08689_),
    .C1(_08666_),
    .X(_00526_));
 sky130_fd_sc_hd__clkbuf_4 _16095_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[3] ),
    .X(_08690_));
 sky130_fd_sc_hd__or2_1 _16096_ (.A(_08690_),
    .B(_08684_),
    .X(_08691_));
 sky130_fd_sc_hd__clkbuf_4 _16097_ (.A(_07617_),
    .X(_08692_));
 sky130_fd_sc_hd__o211a_1 _16098_ (.A1(_08669_),
    .A2(_08681_),
    .B1(_08691_),
    .C1(_08692_),
    .X(_00527_));
 sky130_fd_sc_hd__clkbuf_4 _16099_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[4] ),
    .X(_08693_));
 sky130_fd_sc_hd__or2_1 _16100_ (.A(_08693_),
    .B(_08684_),
    .X(_08694_));
 sky130_fd_sc_hd__o211a_1 _16101_ (.A1(_08671_),
    .A2(_08681_),
    .B1(_08694_),
    .C1(_08692_),
    .X(_00528_));
 sky130_fd_sc_hd__clkbuf_4 _16102_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[5] ),
    .X(_08695_));
 sky130_fd_sc_hd__or2_1 _16103_ (.A(_08695_),
    .B(_08684_),
    .X(_08696_));
 sky130_fd_sc_hd__o211a_1 _16104_ (.A1(_08673_),
    .A2(_08681_),
    .B1(_08696_),
    .C1(_08692_),
    .X(_00529_));
 sky130_fd_sc_hd__buf_2 _16105_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[6] ),
    .X(_08697_));
 sky130_fd_sc_hd__or2_1 _16106_ (.A(_08697_),
    .B(_08684_),
    .X(_08698_));
 sky130_fd_sc_hd__o211a_1 _16107_ (.A1(_08677_),
    .A2(_08681_),
    .B1(_08698_),
    .C1(_08692_),
    .X(_00530_));
 sky130_fd_sc_hd__or2_1 _16108_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[7] ),
    .B(_08684_),
    .X(_08699_));
 sky130_fd_sc_hd__o211a_1 _16109_ (.A1(_08679_),
    .A2(_08681_),
    .B1(_08699_),
    .C1(_08692_),
    .X(_00531_));
 sky130_fd_sc_hd__and3_1 _16110_ (.A(_08683_),
    .B(_08661_),
    .C(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[0] ),
    .X(_08700_));
 sky130_fd_sc_hd__a21oi_1 _16111_ (.A1(_08683_),
    .A2(_08661_),
    .B1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[0] ),
    .Y(_08701_));
 sky130_fd_sc_hd__o21ai_1 _16112_ (.A1(_08700_),
    .A2(_08701_),
    .B1(_08181_),
    .Y(_08702_));
 sky130_fd_sc_hd__o211a_1 _16113_ (.A1(net1068),
    .A2(_08183_),
    .B1(_08702_),
    .C1(_08692_),
    .X(_00532_));
 sky130_fd_sc_hd__a22o_1 _16114_ (.A1(_08664_),
    .A2(_08683_),
    .B1(_08661_),
    .B2(_08686_),
    .X(_08703_));
 sky130_fd_sc_hd__nand4_1 _16115_ (.A(_08686_),
    .B(_08664_),
    .C(_08683_),
    .D(_08661_),
    .Y(_08704_));
 sky130_fd_sc_hd__nand3_1 _16116_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[1] ),
    .B(_08703_),
    .C(_08704_),
    .Y(_08705_));
 sky130_fd_sc_hd__a21o_1 _16117_ (.A1(_08703_),
    .A2(_08704_),
    .B1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[1] ),
    .X(_08706_));
 sky130_fd_sc_hd__a21o_1 _16118_ (.A1(_08705_),
    .A2(_08706_),
    .B1(_08700_),
    .X(_08707_));
 sky130_fd_sc_hd__nand3_1 _16119_ (.A(_08700_),
    .B(_08705_),
    .C(_08706_),
    .Y(_08708_));
 sky130_fd_sc_hd__a21o_1 _16120_ (.A1(_08707_),
    .A2(_08708_),
    .B1(_06682_),
    .X(_08709_));
 sky130_fd_sc_hd__o211a_1 _16121_ (.A1(net1064),
    .A2(_08183_),
    .B1(_08709_),
    .C1(_08692_),
    .X(_00533_));
 sky130_fd_sc_hd__nand2_1 _16122_ (.A(_08688_),
    .B(_08661_),
    .Y(_08710_));
 sky130_fd_sc_hd__a22o_1 _16123_ (.A1(_08686_),
    .A2(_08664_),
    .B1(_08683_),
    .B2(_08667_),
    .X(_08711_));
 sky130_fd_sc_hd__nand4_1 _16124_ (.A(_08667_),
    .B(_08686_),
    .C(_08664_),
    .D(_08683_),
    .Y(_08712_));
 sky130_fd_sc_hd__nand2_1 _16125_ (.A(_08711_),
    .B(_08712_),
    .Y(_08713_));
 sky130_fd_sc_hd__xnor2_1 _16126_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[2] ),
    .B(_08713_),
    .Y(_08714_));
 sky130_fd_sc_hd__nand2_1 _16127_ (.A(_08704_),
    .B(_08705_),
    .Y(_08715_));
 sky130_fd_sc_hd__xnor2_1 _16128_ (.A(_08714_),
    .B(_08715_),
    .Y(_08716_));
 sky130_fd_sc_hd__or2_1 _16129_ (.A(_08710_),
    .B(_08716_),
    .X(_08717_));
 sky130_fd_sc_hd__nand2_1 _16130_ (.A(_08710_),
    .B(_08716_),
    .Y(_08718_));
 sky130_fd_sc_hd__and2_1 _16131_ (.A(_08717_),
    .B(_08718_),
    .X(_08719_));
 sky130_fd_sc_hd__xnor2_1 _16132_ (.A(_08708_),
    .B(_08719_),
    .Y(_08720_));
 sky130_fd_sc_hd__or2_1 _16133_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[2] ),
    .B(_07866_),
    .X(_08721_));
 sky130_fd_sc_hd__o211a_1 _16134_ (.A1(_06848_),
    .A2(_08720_),
    .B1(_08721_),
    .C1(_08692_),
    .X(_00534_));
 sky130_fd_sc_hd__and2b_1 _16135_ (.A_N(_08708_),
    .B(_08719_),
    .X(_08722_));
 sky130_fd_sc_hd__nand2_1 _16136_ (.A(_08714_),
    .B(_08715_),
    .Y(_08723_));
 sky130_fd_sc_hd__a22o_1 _16137_ (.A1(_08688_),
    .A2(_08664_),
    .B1(_08661_),
    .B2(_08690_),
    .X(_08724_));
 sky130_fd_sc_hd__and4_2 _16138_ (.A(_08690_),
    .B(_08688_),
    .C(_08664_),
    .D(_08661_),
    .X(_08725_));
 sky130_fd_sc_hd__inv_2 _16139_ (.A(_08725_),
    .Y(_08726_));
 sky130_fd_sc_hd__nand2_1 _16140_ (.A(_08724_),
    .B(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__a22o_1 _16141_ (.A1(_08667_),
    .A2(_08686_),
    .B1(_08683_),
    .B2(_08669_),
    .X(_08728_));
 sky130_fd_sc_hd__nand4_1 _16142_ (.A(_08669_),
    .B(_08667_),
    .C(_08686_),
    .D(_08683_),
    .Y(_08729_));
 sky130_fd_sc_hd__and3_1 _16143_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[3] ),
    .B(_08728_),
    .C(_08729_),
    .X(_08730_));
 sky130_fd_sc_hd__a21oi_1 _16144_ (.A1(_08728_),
    .A2(_08729_),
    .B1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[3] ),
    .Y(_08731_));
 sky130_fd_sc_hd__or2_2 _16145_ (.A(_08730_),
    .B(_08731_),
    .X(_08732_));
 sky130_fd_sc_hd__a21boi_4 _16146_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[2] ),
    .A2(_08711_),
    .B1_N(_08712_),
    .Y(_08733_));
 sky130_fd_sc_hd__xnor2_2 _16147_ (.A(_08732_),
    .B(_08733_),
    .Y(_08734_));
 sky130_fd_sc_hd__xnor2_1 _16148_ (.A(_08727_),
    .B(_08734_),
    .Y(_08735_));
 sky130_fd_sc_hd__a21o_1 _16149_ (.A1(_08723_),
    .A2(_08717_),
    .B1(_08735_),
    .X(_08736_));
 sky130_fd_sc_hd__nand3_1 _16150_ (.A(_08723_),
    .B(_08717_),
    .C(_08735_),
    .Y(_08737_));
 sky130_fd_sc_hd__nand3_2 _16151_ (.A(_08722_),
    .B(_08736_),
    .C(_08737_),
    .Y(_08738_));
 sky130_fd_sc_hd__a21o_1 _16152_ (.A1(_08736_),
    .A2(_08737_),
    .B1(_08722_),
    .X(_08739_));
 sky130_fd_sc_hd__and2_1 _16153_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[3] ),
    .B(_05730_),
    .X(_08740_));
 sky130_fd_sc_hd__a31o_1 _16154_ (.A1(_05887_),
    .A2(_08738_),
    .A3(_08739_),
    .B1(_08740_),
    .X(_08741_));
 sky130_fd_sc_hd__and2_1 _16155_ (.A(_08197_),
    .B(_08741_),
    .X(_08742_));
 sky130_fd_sc_hd__clkbuf_1 _16156_ (.A(_08742_),
    .X(_00535_));
 sky130_fd_sc_hd__a22o_1 _16157_ (.A1(\top_inst.grid_inst.data_path_wires[8][3] ),
    .A2(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[1] ),
    .B1(_08682_),
    .B2(\top_inst.grid_inst.data_path_wires[8][4] ),
    .X(_08743_));
 sky130_fd_sc_hd__nand4_1 _16158_ (.A(_08671_),
    .B(_08669_),
    .C(_08686_),
    .D(_08682_),
    .Y(_08744_));
 sky130_fd_sc_hd__nand2_1 _16159_ (.A(_08743_),
    .B(_08744_),
    .Y(_08745_));
 sky130_fd_sc_hd__xor2_2 _16160_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[4] ),
    .B(_08745_),
    .X(_08746_));
 sky130_fd_sc_hd__xnor2_2 _16161_ (.A(_08725_),
    .B(_08746_),
    .Y(_08747_));
 sky130_fd_sc_hd__a21bo_1 _16162_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[3] ),
    .A2(_08728_),
    .B1_N(_08729_),
    .X(_08748_));
 sky130_fd_sc_hd__xnor2_2 _16163_ (.A(_08747_),
    .B(_08748_),
    .Y(_08749_));
 sky130_fd_sc_hd__nand2_1 _16164_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[2] ),
    .B(_08667_),
    .Y(_08750_));
 sky130_fd_sc_hd__nand4_1 _16165_ (.A(_08693_),
    .B(_08690_),
    .C(\top_inst.grid_inst.data_path_wires[8][1] ),
    .D(\top_inst.grid_inst.data_path_wires[8][0] ),
    .Y(_08751_));
 sky130_fd_sc_hd__a22o_1 _16166_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[3] ),
    .A2(\top_inst.grid_inst.data_path_wires[8][1] ),
    .B1(\top_inst.grid_inst.data_path_wires[8][0] ),
    .B2(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[4] ),
    .X(_08752_));
 sky130_fd_sc_hd__nand2_1 _16167_ (.A(_08751_),
    .B(_08752_),
    .Y(_08753_));
 sky130_fd_sc_hd__xor2_2 _16168_ (.A(_08750_),
    .B(_08753_),
    .X(_08754_));
 sky130_fd_sc_hd__xnor2_2 _16169_ (.A(_08749_),
    .B(_08754_),
    .Y(_08755_));
 sky130_fd_sc_hd__inv_2 _16170_ (.A(_08724_),
    .Y(_08756_));
 sky130_fd_sc_hd__o32ai_4 _16171_ (.A1(_08756_),
    .A2(_08725_),
    .A3(_08734_),
    .B1(_08733_),
    .B2(_08732_),
    .Y(_08757_));
 sky130_fd_sc_hd__xnor2_2 _16172_ (.A(_08755_),
    .B(_08757_),
    .Y(_08758_));
 sky130_fd_sc_hd__nand2_1 _16173_ (.A(_08736_),
    .B(_08738_),
    .Y(_08759_));
 sky130_fd_sc_hd__nor2_1 _16174_ (.A(_08758_),
    .B(_08759_),
    .Y(_08760_));
 sky130_fd_sc_hd__a21o_1 _16175_ (.A1(_08758_),
    .A2(_08759_),
    .B1(_07057_),
    .X(_08761_));
 sky130_fd_sc_hd__o221a_1 _16176_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[4] ),
    .A2(_07048_),
    .B1(_08760_),
    .B2(_08761_),
    .C1(_07708_),
    .X(_00536_));
 sky130_fd_sc_hd__nor2_1 _16177_ (.A(_08738_),
    .B(_08758_),
    .Y(_08762_));
 sky130_fd_sc_hd__and2b_1 _16178_ (.A_N(_08749_),
    .B(_08754_),
    .X(_08763_));
 sky130_fd_sc_hd__nand2_1 _16179_ (.A(_08695_),
    .B(_08661_),
    .Y(_08764_));
 sky130_fd_sc_hd__a22o_1 _16180_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[3] ),
    .A2(\top_inst.grid_inst.data_path_wires[8][2] ),
    .B1(\top_inst.grid_inst.data_path_wires[8][1] ),
    .B2(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[4] ),
    .X(_08765_));
 sky130_fd_sc_hd__nand4_1 _16181_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[3] ),
    .C(_08667_),
    .D(\top_inst.grid_inst.data_path_wires[8][1] ),
    .Y(_08766_));
 sky130_fd_sc_hd__nand2_1 _16182_ (.A(_08765_),
    .B(_08766_),
    .Y(_08767_));
 sky130_fd_sc_hd__nand2_1 _16183_ (.A(_08669_),
    .B(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[2] ),
    .Y(_08768_));
 sky130_fd_sc_hd__xor2_1 _16184_ (.A(_08767_),
    .B(_08768_),
    .X(_08769_));
 sky130_fd_sc_hd__xnor2_1 _16185_ (.A(_08764_),
    .B(_08769_),
    .Y(_08770_));
 sky130_fd_sc_hd__a21boi_2 _16186_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[4] ),
    .A2(_08743_),
    .B1_N(_08744_),
    .Y(_08771_));
 sky130_fd_sc_hd__o21ai_1 _16187_ (.A1(_08750_),
    .A2(_08753_),
    .B1(_08751_),
    .Y(_08772_));
 sky130_fd_sc_hd__a22o_1 _16188_ (.A1(\top_inst.grid_inst.data_path_wires[8][4] ),
    .A2(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[1] ),
    .B1(_08682_),
    .B2(\top_inst.grid_inst.data_path_wires[8][5] ),
    .X(_08773_));
 sky130_fd_sc_hd__nand4_1 _16189_ (.A(_08673_),
    .B(\top_inst.grid_inst.data_path_wires[8][4] ),
    .C(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[1] ),
    .D(_08682_),
    .Y(_08774_));
 sky130_fd_sc_hd__nand2_1 _16190_ (.A(_08773_),
    .B(_08774_),
    .Y(_08775_));
 sky130_fd_sc_hd__xor2_2 _16191_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[5] ),
    .B(_08775_),
    .X(_08776_));
 sky130_fd_sc_hd__xnor2_1 _16192_ (.A(_08772_),
    .B(_08776_),
    .Y(_08777_));
 sky130_fd_sc_hd__xnor2_1 _16193_ (.A(_08771_),
    .B(_08777_),
    .Y(_08778_));
 sky130_fd_sc_hd__xor2_1 _16194_ (.A(_08770_),
    .B(_08778_),
    .X(_08779_));
 sky130_fd_sc_hd__xor2_1 _16195_ (.A(_08763_),
    .B(_08779_),
    .X(_08780_));
 sky130_fd_sc_hd__nor2_1 _16196_ (.A(_08726_),
    .B(_08746_),
    .Y(_08781_));
 sky130_fd_sc_hd__a21o_1 _16197_ (.A1(_08747_),
    .A2(_08748_),
    .B1(_08781_),
    .X(_08782_));
 sky130_fd_sc_hd__xnor2_1 _16198_ (.A(_08780_),
    .B(_08782_),
    .Y(_08783_));
 sky130_fd_sc_hd__nand2_1 _16199_ (.A(_08755_),
    .B(_08757_),
    .Y(_08784_));
 sky130_fd_sc_hd__o21ai_1 _16200_ (.A1(_08736_),
    .A2(_08758_),
    .B1(_08784_),
    .Y(_08785_));
 sky130_fd_sc_hd__xnor2_1 _16201_ (.A(_08783_),
    .B(_08785_),
    .Y(_08786_));
 sky130_fd_sc_hd__nand2_1 _16202_ (.A(_08762_),
    .B(_08786_),
    .Y(_08787_));
 sky130_fd_sc_hd__o21a_1 _16203_ (.A1(_08762_),
    .A2(_08786_),
    .B1(_08265_),
    .X(_08788_));
 sky130_fd_sc_hd__a22o_1 _16204_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[5] ),
    .A2(_08066_),
    .B1(_08787_),
    .B2(_08788_),
    .X(_08789_));
 sky130_fd_sc_hd__and2_1 _16205_ (.A(_08197_),
    .B(_08789_),
    .X(_08790_));
 sky130_fd_sc_hd__clkbuf_1 _16206_ (.A(_08790_),
    .X(_00537_));
 sky130_fd_sc_hd__nor2_1 _16207_ (.A(_08784_),
    .B(_08783_),
    .Y(_08791_));
 sky130_fd_sc_hd__nand2_1 _16208_ (.A(_08763_),
    .B(_08779_),
    .Y(_08792_));
 sky130_fd_sc_hd__nand2_1 _16209_ (.A(_08780_),
    .B(_08782_),
    .Y(_08793_));
 sky130_fd_sc_hd__or2b_1 _16210_ (.A(_08776_),
    .B_N(_08772_),
    .X(_08794_));
 sky130_fd_sc_hd__or2b_1 _16211_ (.A(_08771_),
    .B_N(_08777_),
    .X(_08795_));
 sky130_fd_sc_hd__or2b_1 _16212_ (.A(_08764_),
    .B_N(_08769_),
    .X(_08796_));
 sky130_fd_sc_hd__a22o_1 _16213_ (.A1(_08695_),
    .A2(_08664_),
    .B1(\top_inst.grid_inst.data_path_wires[8][0] ),
    .B2(_08697_),
    .X(_08797_));
 sky130_fd_sc_hd__nand4_2 _16214_ (.A(_08697_),
    .B(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[5] ),
    .C(_08664_),
    .D(\top_inst.grid_inst.data_path_wires[8][0] ),
    .Y(_08798_));
 sky130_fd_sc_hd__nand2_1 _16215_ (.A(_08797_),
    .B(_08798_),
    .Y(_08799_));
 sky130_fd_sc_hd__a22o_1 _16216_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[3] ),
    .A2(\top_inst.grid_inst.data_path_wires[8][3] ),
    .B1(_08667_),
    .B2(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[4] ),
    .X(_08800_));
 sky130_fd_sc_hd__nand4_2 _16217_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[3] ),
    .C(\top_inst.grid_inst.data_path_wires[8][3] ),
    .D(_08667_),
    .Y(_08801_));
 sky130_fd_sc_hd__a22o_1 _16218_ (.A1(_08671_),
    .A2(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[2] ),
    .B1(_08800_),
    .B2(_08801_),
    .X(_08802_));
 sky130_fd_sc_hd__nand4_2 _16219_ (.A(_08671_),
    .B(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[2] ),
    .C(_08800_),
    .D(_08801_),
    .Y(_08803_));
 sky130_fd_sc_hd__nand2_1 _16220_ (.A(_08802_),
    .B(_08803_),
    .Y(_08804_));
 sky130_fd_sc_hd__xnor2_1 _16221_ (.A(_08799_),
    .B(_08804_),
    .Y(_08805_));
 sky130_fd_sc_hd__xor2_1 _16222_ (.A(_08796_),
    .B(_08805_),
    .X(_08806_));
 sky130_fd_sc_hd__a21boi_2 _16223_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[5] ),
    .A2(_08773_),
    .B1_N(_08774_),
    .Y(_08807_));
 sky130_fd_sc_hd__o21a_1 _16224_ (.A1(_08767_),
    .A2(_08768_),
    .B1(_08766_),
    .X(_08808_));
 sky130_fd_sc_hd__a22o_1 _16225_ (.A1(\top_inst.grid_inst.data_path_wires[8][5] ),
    .A2(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[1] ),
    .B1(_08682_),
    .B2(_08676_),
    .X(_08809_));
 sky130_fd_sc_hd__nand4_1 _16226_ (.A(_08676_),
    .B(\top_inst.grid_inst.data_path_wires[8][5] ),
    .C(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[1] ),
    .D(_08682_),
    .Y(_08810_));
 sky130_fd_sc_hd__nand2_1 _16227_ (.A(_08809_),
    .B(_08810_),
    .Y(_08811_));
 sky130_fd_sc_hd__xor2_2 _16228_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[6] ),
    .B(_08811_),
    .X(_08812_));
 sky130_fd_sc_hd__xor2_1 _16229_ (.A(_08808_),
    .B(_08812_),
    .X(_08813_));
 sky130_fd_sc_hd__xnor2_1 _16230_ (.A(_08807_),
    .B(_08813_),
    .Y(_08814_));
 sky130_fd_sc_hd__nand2_1 _16231_ (.A(_08806_),
    .B(_08814_),
    .Y(_08815_));
 sky130_fd_sc_hd__or2_1 _16232_ (.A(_08806_),
    .B(_08814_),
    .X(_08816_));
 sky130_fd_sc_hd__and2_1 _16233_ (.A(_08770_),
    .B(_08778_),
    .X(_08817_));
 sky130_fd_sc_hd__a21oi_1 _16234_ (.A1(_08815_),
    .A2(_08816_),
    .B1(_08817_),
    .Y(_08818_));
 sky130_fd_sc_hd__and3_1 _16235_ (.A(_08817_),
    .B(_08815_),
    .C(_08816_),
    .X(_08819_));
 sky130_fd_sc_hd__a211oi_2 _16236_ (.A1(_08794_),
    .A2(_08795_),
    .B1(_08818_),
    .C1(_08819_),
    .Y(_08820_));
 sky130_fd_sc_hd__o211a_1 _16237_ (.A1(_08818_),
    .A2(_08819_),
    .B1(_08794_),
    .C1(_08795_),
    .X(_08821_));
 sky130_fd_sc_hd__a211o_1 _16238_ (.A1(_08792_),
    .A2(_08793_),
    .B1(_08820_),
    .C1(_08821_),
    .X(_08822_));
 sky130_fd_sc_hd__o211ai_1 _16239_ (.A1(_08820_),
    .A2(_08821_),
    .B1(_08792_),
    .C1(_08793_),
    .Y(_08823_));
 sky130_fd_sc_hd__and3_1 _16240_ (.A(_08791_),
    .B(_08822_),
    .C(_08823_),
    .X(_08824_));
 sky130_fd_sc_hd__a21oi_1 _16241_ (.A1(_08822_),
    .A2(_08823_),
    .B1(_08791_),
    .Y(_08825_));
 sky130_fd_sc_hd__nor2_1 _16242_ (.A(_08824_),
    .B(_08825_),
    .Y(_08826_));
 sky130_fd_sc_hd__o31a_1 _16243_ (.A1(_08736_),
    .A2(_08758_),
    .A3(_08783_),
    .B1(_08787_),
    .X(_08827_));
 sky130_fd_sc_hd__xnor2_1 _16244_ (.A(_08826_),
    .B(_08827_),
    .Y(_08828_));
 sky130_fd_sc_hd__mux2_1 _16245_ (.A0(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[6] ),
    .A1(_08828_),
    .S(_08307_),
    .X(_08829_));
 sky130_fd_sc_hd__and2_1 _16246_ (.A(_08197_),
    .B(_08829_),
    .X(_08830_));
 sky130_fd_sc_hd__clkbuf_1 _16247_ (.A(_08830_),
    .X(_00538_));
 sky130_fd_sc_hd__clkbuf_4 _16248_ (.A(_04873_),
    .X(_08831_));
 sky130_fd_sc_hd__nor2_1 _16249_ (.A(_08799_),
    .B(_08804_),
    .Y(_08832_));
 sky130_fd_sc_hd__nand2_1 _16250_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[6] ),
    .B(\top_inst.grid_inst.data_path_wires[8][1] ),
    .Y(_08833_));
 sky130_fd_sc_hd__or2b_1 _16251_ (.A(\top_inst.grid_inst.data_path_wires[8][0] ),
    .B_N(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[7] ),
    .X(_08834_));
 sky130_fd_sc_hd__xnor2_1 _16252_ (.A(_08833_),
    .B(_08834_),
    .Y(_08835_));
 sky130_fd_sc_hd__nand2_1 _16253_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[5] ),
    .B(\top_inst.grid_inst.data_path_wires[8][2] ),
    .Y(_08836_));
 sky130_fd_sc_hd__xnor2_1 _16254_ (.A(_08835_),
    .B(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__xor2_1 _16255_ (.A(_08798_),
    .B(_08837_),
    .X(_08838_));
 sky130_fd_sc_hd__a22o_1 _16256_ (.A1(\top_inst.grid_inst.data_path_wires[8][4] ),
    .A2(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[3] ),
    .B1(\top_inst.grid_inst.data_path_wires[8][3] ),
    .B2(_08693_),
    .X(_08839_));
 sky130_fd_sc_hd__nand4_2 _16257_ (.A(_08693_),
    .B(\top_inst.grid_inst.data_path_wires[8][4] ),
    .C(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[3] ),
    .D(_08669_),
    .Y(_08840_));
 sky130_fd_sc_hd__a22o_1 _16258_ (.A1(_08673_),
    .A2(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[2] ),
    .B1(_08839_),
    .B2(_08840_),
    .X(_08841_));
 sky130_fd_sc_hd__nand4_2 _16259_ (.A(_08673_),
    .B(_08688_),
    .C(_08839_),
    .D(_08840_),
    .Y(_08842_));
 sky130_fd_sc_hd__nand2_1 _16260_ (.A(_08841_),
    .B(_08842_),
    .Y(_08843_));
 sky130_fd_sc_hd__xnor2_1 _16261_ (.A(_08838_),
    .B(_08843_),
    .Y(_08844_));
 sky130_fd_sc_hd__xnor2_1 _16262_ (.A(_08832_),
    .B(_08844_),
    .Y(_08845_));
 sky130_fd_sc_hd__a21bo_1 _16263_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[6] ),
    .A2(_08809_),
    .B1_N(_08810_),
    .X(_08846_));
 sky130_fd_sc_hd__a22o_1 _16264_ (.A1(_08676_),
    .A2(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[1] ),
    .B1(_08682_),
    .B2(\top_inst.grid_inst.data_path_wires[8][7] ),
    .X(_08847_));
 sky130_fd_sc_hd__nand4_1 _16265_ (.A(\top_inst.grid_inst.data_path_wires[8][7] ),
    .B(_08676_),
    .C(_08686_),
    .D(_08682_),
    .Y(_08848_));
 sky130_fd_sc_hd__and3_1 _16266_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[7] ),
    .B(_08847_),
    .C(_08848_),
    .X(_08849_));
 sky130_fd_sc_hd__a21oi_1 _16267_ (.A1(_08847_),
    .A2(_08848_),
    .B1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[7] ),
    .Y(_08850_));
 sky130_fd_sc_hd__a211oi_1 _16268_ (.A1(_08801_),
    .A2(_08803_),
    .B1(_08849_),
    .C1(_08850_),
    .Y(_08851_));
 sky130_fd_sc_hd__o211a_1 _16269_ (.A1(_08849_),
    .A2(_08850_),
    .B1(_08801_),
    .C1(_08803_),
    .X(_08852_));
 sky130_fd_sc_hd__nor2_1 _16270_ (.A(_08851_),
    .B(_08852_),
    .Y(_08853_));
 sky130_fd_sc_hd__xnor2_1 _16271_ (.A(_08846_),
    .B(_08853_),
    .Y(_08854_));
 sky130_fd_sc_hd__xor2_1 _16272_ (.A(_08845_),
    .B(_08854_),
    .X(_08855_));
 sky130_fd_sc_hd__o21ai_1 _16273_ (.A1(_08796_),
    .A2(_08805_),
    .B1(_08815_),
    .Y(_08856_));
 sky130_fd_sc_hd__xnor2_1 _16274_ (.A(_08855_),
    .B(_08856_),
    .Y(_08857_));
 sky130_fd_sc_hd__or2b_1 _16275_ (.A(_08807_),
    .B_N(_08813_),
    .X(_08858_));
 sky130_fd_sc_hd__o21ai_1 _16276_ (.A1(_08808_),
    .A2(_08812_),
    .B1(_08858_),
    .Y(_08859_));
 sky130_fd_sc_hd__xnor2_1 _16277_ (.A(_08857_),
    .B(_08859_),
    .Y(_08860_));
 sky130_fd_sc_hd__nor2_1 _16278_ (.A(_08819_),
    .B(_08820_),
    .Y(_08861_));
 sky130_fd_sc_hd__xnor2_1 _16279_ (.A(_08860_),
    .B(_08861_),
    .Y(_08862_));
 sky130_fd_sc_hd__xnor2_1 _16280_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[7] ),
    .B(_08862_),
    .Y(_08863_));
 sky130_fd_sc_hd__xor2_1 _16281_ (.A(_08822_),
    .B(_08863_),
    .X(_08864_));
 sky130_fd_sc_hd__o21bai_1 _16282_ (.A1(_08825_),
    .A2(_08827_),
    .B1_N(_08824_),
    .Y(_08865_));
 sky130_fd_sc_hd__nor2_1 _16283_ (.A(_08864_),
    .B(_08865_),
    .Y(_08866_));
 sky130_fd_sc_hd__a21o_1 _16284_ (.A1(_08864_),
    .A2(_08865_),
    .B1(_05353_),
    .X(_08867_));
 sky130_fd_sc_hd__a2bb2o_1 _16285_ (.A1_N(_08866_),
    .A2_N(_08867_),
    .B1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[7] ),
    .B2(_07816_),
    .X(_08868_));
 sky130_fd_sc_hd__and2_1 _16286_ (.A(_08831_),
    .B(_08868_),
    .X(_08869_));
 sky130_fd_sc_hd__clkbuf_1 _16287_ (.A(_08869_),
    .X(_00539_));
 sky130_fd_sc_hd__buf_4 _16288_ (.A(_05732_),
    .X(_08870_));
 sky130_fd_sc_hd__nor2_1 _16289_ (.A(_08822_),
    .B(_08863_),
    .Y(_08871_));
 sky130_fd_sc_hd__a21o_1 _16290_ (.A1(_08864_),
    .A2(_08865_),
    .B1(_08871_),
    .X(_08872_));
 sky130_fd_sc_hd__or2b_1 _16291_ (.A(_08861_),
    .B_N(_08860_),
    .X(_08873_));
 sky130_fd_sc_hd__nand2_1 _16292_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[7] ),
    .B(_08862_),
    .Y(_08874_));
 sky130_fd_sc_hd__and4b_1 _16293_ (.A_N(\top_inst.grid_inst.data_path_wires[8][1] ),
    .B(\top_inst.grid_inst.data_path_wires[8][2] ),
    .C(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[6] ),
    .D(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[7] ),
    .X(_08875_));
 sky130_fd_sc_hd__inv_2 _16294_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[7] ),
    .Y(_08876_));
 sky130_fd_sc_hd__o2bb2a_1 _16295_ (.A1_N(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[6] ),
    .A2_N(\top_inst.grid_inst.data_path_wires[8][2] ),
    .B1(\top_inst.grid_inst.data_path_wires[8][1] ),
    .B2(_08876_),
    .X(_08877_));
 sky130_fd_sc_hd__nor2_2 _16296_ (.A(_08875_),
    .B(_08877_),
    .Y(_08878_));
 sky130_fd_sc_hd__nand2_2 _16297_ (.A(_08695_),
    .B(_08669_),
    .Y(_08879_));
 sky130_fd_sc_hd__xnor2_4 _16298_ (.A(_08878_),
    .B(_08879_),
    .Y(_08880_));
 sky130_fd_sc_hd__nor2_1 _16299_ (.A(_08835_),
    .B(_08836_),
    .Y(_08881_));
 sky130_fd_sc_hd__o21ba_1 _16300_ (.A1(_08833_),
    .A2(_08834_),
    .B1_N(_08881_),
    .X(_08882_));
 sky130_fd_sc_hd__xnor2_2 _16301_ (.A(_08880_),
    .B(_08882_),
    .Y(_08883_));
 sky130_fd_sc_hd__a22o_1 _16302_ (.A1(_08693_),
    .A2(_08671_),
    .B1(_08690_),
    .B2(_08673_),
    .X(_08884_));
 sky130_fd_sc_hd__nand4_4 _16303_ (.A(_08673_),
    .B(_08693_),
    .C(_08671_),
    .D(_08690_),
    .Y(_08885_));
 sky130_fd_sc_hd__a22o_1 _16304_ (.A1(_08677_),
    .A2(_08688_),
    .B1(_08884_),
    .B2(_08885_),
    .X(_08886_));
 sky130_fd_sc_hd__nand4_4 _16305_ (.A(_08677_),
    .B(_08688_),
    .C(_08884_),
    .D(_08885_),
    .Y(_08887_));
 sky130_fd_sc_hd__nand2_1 _16306_ (.A(_08886_),
    .B(_08887_),
    .Y(_08888_));
 sky130_fd_sc_hd__xnor2_1 _16307_ (.A(_08883_),
    .B(_08888_),
    .Y(_08889_));
 sky130_fd_sc_hd__and3_1 _16308_ (.A(_08838_),
    .B(_08841_),
    .C(_08842_),
    .X(_08890_));
 sky130_fd_sc_hd__o21ba_1 _16309_ (.A1(_08798_),
    .A2(_08837_),
    .B1_N(_08890_),
    .X(_08891_));
 sky130_fd_sc_hd__xnor2_1 _16310_ (.A(_08889_),
    .B(_08891_),
    .Y(_08892_));
 sky130_fd_sc_hd__and4_1 _16311_ (.A(_08679_),
    .B(_08677_),
    .C(_08686_),
    .D(_08683_),
    .X(_08893_));
 sky130_fd_sc_hd__o21ai_2 _16312_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[1] ),
    .A2(_08682_),
    .B1(\top_inst.grid_inst.data_path_wires[8][7] ),
    .Y(_08894_));
 sky130_fd_sc_hd__and3_1 _16313_ (.A(\top_inst.grid_inst.data_path_wires[8][7] ),
    .B(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[1] ),
    .C(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[0] ),
    .X(_08895_));
 sky130_fd_sc_hd__buf_4 _16314_ (.A(_08895_),
    .X(_08896_));
 sky130_fd_sc_hd__nor2_4 _16315_ (.A(_08894_),
    .B(_08896_),
    .Y(_08897_));
 sky130_fd_sc_hd__xnor2_1 _16316_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[8] ),
    .B(_08897_),
    .Y(_08898_));
 sky130_fd_sc_hd__a21oi_1 _16317_ (.A1(_08840_),
    .A2(_08842_),
    .B1(_08898_),
    .Y(_08899_));
 sky130_fd_sc_hd__and3_1 _16318_ (.A(_08840_),
    .B(_08842_),
    .C(_08898_),
    .X(_08900_));
 sky130_fd_sc_hd__nor2_1 _16319_ (.A(_08899_),
    .B(_08900_),
    .Y(_08901_));
 sky130_fd_sc_hd__o21a_1 _16320_ (.A1(_08893_),
    .A2(_08849_),
    .B1(_08901_),
    .X(_08902_));
 sky130_fd_sc_hd__nor3_1 _16321_ (.A(_08893_),
    .B(_08849_),
    .C(_08901_),
    .Y(_08903_));
 sky130_fd_sc_hd__nor2_1 _16322_ (.A(_08902_),
    .B(_08903_),
    .Y(_08904_));
 sky130_fd_sc_hd__xnor2_1 _16323_ (.A(_08892_),
    .B(_08904_),
    .Y(_08905_));
 sky130_fd_sc_hd__nand2_1 _16324_ (.A(_08832_),
    .B(_08844_),
    .Y(_08906_));
 sky130_fd_sc_hd__o21a_1 _16325_ (.A1(_08845_),
    .A2(_08854_),
    .B1(_08906_),
    .X(_08907_));
 sky130_fd_sc_hd__xnor2_1 _16326_ (.A(_08905_),
    .B(_08907_),
    .Y(_08908_));
 sky130_fd_sc_hd__a21oi_1 _16327_ (.A1(_08846_),
    .A2(_08853_),
    .B1(_08851_),
    .Y(_08909_));
 sky130_fd_sc_hd__xnor2_1 _16328_ (.A(_08908_),
    .B(_08909_),
    .Y(_08910_));
 sky130_fd_sc_hd__and2b_1 _16329_ (.A_N(_08857_),
    .B(_08859_),
    .X(_08911_));
 sky130_fd_sc_hd__a21oi_1 _16330_ (.A1(_08855_),
    .A2(_08856_),
    .B1(_08911_),
    .Y(_08912_));
 sky130_fd_sc_hd__xnor2_1 _16331_ (.A(_08910_),
    .B(_08912_),
    .Y(_08913_));
 sky130_fd_sc_hd__a21o_1 _16332_ (.A1(_08873_),
    .A2(_08874_),
    .B1(_08913_),
    .X(_08914_));
 sky130_fd_sc_hd__nand3_1 _16333_ (.A(_08873_),
    .B(_08874_),
    .C(_08913_),
    .Y(_08915_));
 sky130_fd_sc_hd__and2_1 _16334_ (.A(_08914_),
    .B(_08915_),
    .X(_08916_));
 sky130_fd_sc_hd__xor2_1 _16335_ (.A(_08872_),
    .B(_08916_),
    .X(_08917_));
 sky130_fd_sc_hd__or2_1 _16336_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[8] ),
    .B(_07866_),
    .X(_08918_));
 sky130_fd_sc_hd__o211a_1 _16337_ (.A1(_08870_),
    .A2(_08917_),
    .B1(_08918_),
    .C1(_08692_),
    .X(_00540_));
 sky130_fd_sc_hd__a21bo_1 _16338_ (.A1(_08872_),
    .A2(_08916_),
    .B1_N(_08914_),
    .X(_08919_));
 sky130_fd_sc_hd__or2_1 _16339_ (.A(_08910_),
    .B(_08912_),
    .X(_08920_));
 sky130_fd_sc_hd__and4b_1 _16340_ (.A_N(\top_inst.grid_inst.data_path_wires[8][2] ),
    .B(\top_inst.grid_inst.data_path_wires[8][3] ),
    .C(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[6] ),
    .D(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[7] ),
    .X(_08921_));
 sky130_fd_sc_hd__o2bb2a_1 _16341_ (.A1_N(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[6] ),
    .A2_N(\top_inst.grid_inst.data_path_wires[8][3] ),
    .B1(\top_inst.grid_inst.data_path_wires[8][2] ),
    .B2(_08876_),
    .X(_08922_));
 sky130_fd_sc_hd__nor2_1 _16342_ (.A(_08921_),
    .B(_08922_),
    .Y(_08923_));
 sky130_fd_sc_hd__nand2_1 _16343_ (.A(_08695_),
    .B(_08671_),
    .Y(_08924_));
 sky130_fd_sc_hd__xnor2_1 _16344_ (.A(_08923_),
    .B(_08924_),
    .Y(_08925_));
 sky130_fd_sc_hd__o21ba_1 _16345_ (.A1(_08877_),
    .A2(_08879_),
    .B1_N(_08875_),
    .X(_08926_));
 sky130_fd_sc_hd__xor2_1 _16346_ (.A(_08925_),
    .B(_08926_),
    .X(_08927_));
 sky130_fd_sc_hd__a22o_1 _16347_ (.A1(_08673_),
    .A2(_08693_),
    .B1(_08690_),
    .B2(_08676_),
    .X(_08928_));
 sky130_fd_sc_hd__and4_1 _16348_ (.A(\top_inst.grid_inst.data_path_wires[8][6] ),
    .B(\top_inst.grid_inst.data_path_wires[8][5] ),
    .C(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[3] ),
    .X(_08929_));
 sky130_fd_sc_hd__inv_2 _16349_ (.A(_08929_),
    .Y(_08930_));
 sky130_fd_sc_hd__and2_1 _16350_ (.A(_08928_),
    .B(_08930_),
    .X(_08931_));
 sky130_fd_sc_hd__nand2_4 _16351_ (.A(\top_inst.grid_inst.data_path_wires[8][7] ),
    .B(_08688_),
    .Y(_08932_));
 sky130_fd_sc_hd__xor2_1 _16352_ (.A(_08931_),
    .B(_08932_),
    .X(_08933_));
 sky130_fd_sc_hd__xor2_1 _16353_ (.A(_08927_),
    .B(_08933_),
    .X(_08934_));
 sky130_fd_sc_hd__inv_2 _16354_ (.A(_08882_),
    .Y(_08935_));
 sky130_fd_sc_hd__a32oi_4 _16355_ (.A1(_08883_),
    .A2(_08886_),
    .A3(_08887_),
    .B1(_08935_),
    .B2(_08880_),
    .Y(_08936_));
 sky130_fd_sc_hd__xnor2_1 _16356_ (.A(_08934_),
    .B(_08936_),
    .Y(_08937_));
 sky130_fd_sc_hd__a21o_1 _16357_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[8] ),
    .A2(_08897_),
    .B1(_08896_),
    .X(_08938_));
 sky130_fd_sc_hd__xnor2_1 _16358_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[9] ),
    .B(_08897_),
    .Y(_08939_));
 sky130_fd_sc_hd__a21oi_1 _16359_ (.A1(_08885_),
    .A2(_08887_),
    .B1(_08939_),
    .Y(_08940_));
 sky130_fd_sc_hd__and3_1 _16360_ (.A(_08885_),
    .B(_08887_),
    .C(_08939_),
    .X(_08941_));
 sky130_fd_sc_hd__nor2_1 _16361_ (.A(_08940_),
    .B(_08941_),
    .Y(_08942_));
 sky130_fd_sc_hd__xor2_1 _16362_ (.A(_08938_),
    .B(_08942_),
    .X(_08943_));
 sky130_fd_sc_hd__xnor2_1 _16363_ (.A(_08937_),
    .B(_08943_),
    .Y(_08944_));
 sky130_fd_sc_hd__and2b_1 _16364_ (.A_N(_08891_),
    .B(_08889_),
    .X(_08945_));
 sky130_fd_sc_hd__a21oi_1 _16365_ (.A1(_08892_),
    .A2(_08904_),
    .B1(_08945_),
    .Y(_08946_));
 sky130_fd_sc_hd__xnor2_1 _16366_ (.A(_08944_),
    .B(_08946_),
    .Y(_08947_));
 sky130_fd_sc_hd__nor2_1 _16367_ (.A(_08899_),
    .B(_08902_),
    .Y(_08948_));
 sky130_fd_sc_hd__xnor2_1 _16368_ (.A(_08947_),
    .B(_08948_),
    .Y(_08949_));
 sky130_fd_sc_hd__or2_1 _16369_ (.A(_08905_),
    .B(_08907_),
    .X(_08950_));
 sky130_fd_sc_hd__o21a_1 _16370_ (.A1(_08908_),
    .A2(_08909_),
    .B1(_08950_),
    .X(_08951_));
 sky130_fd_sc_hd__nor2_1 _16371_ (.A(_08949_),
    .B(_08951_),
    .Y(_08952_));
 sky130_fd_sc_hd__and2_1 _16372_ (.A(_08949_),
    .B(_08951_),
    .X(_08953_));
 sky130_fd_sc_hd__or2_1 _16373_ (.A(_08952_),
    .B(_08953_),
    .X(_08954_));
 sky130_fd_sc_hd__xor2_1 _16374_ (.A(_08920_),
    .B(_08954_),
    .X(_08955_));
 sky130_fd_sc_hd__xor2_1 _16375_ (.A(_08919_),
    .B(_08955_),
    .X(_08956_));
 sky130_fd_sc_hd__or2_1 _16376_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[9] ),
    .B(_07866_),
    .X(_08957_));
 sky130_fd_sc_hd__o211a_1 _16377_ (.A1(_08870_),
    .A2(_08956_),
    .B1(_08957_),
    .C1(_08692_),
    .X(_00541_));
 sky130_fd_sc_hd__or2b_1 _16378_ (.A(_08926_),
    .B_N(_08925_),
    .X(_08958_));
 sky130_fd_sc_hd__o21a_1 _16379_ (.A1(_08927_),
    .A2(_08933_),
    .B1(_08958_),
    .X(_08959_));
 sky130_fd_sc_hd__and4b_1 _16380_ (.A_N(_08669_),
    .B(_08671_),
    .C(_08697_),
    .D(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[7] ),
    .X(_08960_));
 sky130_fd_sc_hd__o2bb2a_1 _16381_ (.A1_N(_08697_),
    .A2_N(_08671_),
    .B1(_08669_),
    .B2(_08876_),
    .X(_08961_));
 sky130_fd_sc_hd__nor2_1 _16382_ (.A(_08960_),
    .B(_08961_),
    .Y(_08962_));
 sky130_fd_sc_hd__nand2_1 _16383_ (.A(_08695_),
    .B(_08673_),
    .Y(_08963_));
 sky130_fd_sc_hd__xnor2_1 _16384_ (.A(_08962_),
    .B(_08963_),
    .Y(_08964_));
 sky130_fd_sc_hd__o21ba_1 _16385_ (.A1(_08922_),
    .A2(_08924_),
    .B1_N(_08921_),
    .X(_08965_));
 sky130_fd_sc_hd__xnor2_1 _16386_ (.A(_08964_),
    .B(_08965_),
    .Y(_08966_));
 sky130_fd_sc_hd__and3_1 _16387_ (.A(\top_inst.grid_inst.data_path_wires[8][7] ),
    .B(_08693_),
    .C(_08690_),
    .X(_08967_));
 sky130_fd_sc_hd__a22o_1 _16388_ (.A1(_08676_),
    .A2(_08693_),
    .B1(_08690_),
    .B2(\top_inst.grid_inst.data_path_wires[8][7] ),
    .X(_08968_));
 sky130_fd_sc_hd__a21bo_1 _16389_ (.A1(_08677_),
    .A2(_08967_),
    .B1_N(_08968_),
    .X(_08969_));
 sky130_fd_sc_hd__xor2_1 _16390_ (.A(_08932_),
    .B(_08969_),
    .X(_08970_));
 sky130_fd_sc_hd__xor2_1 _16391_ (.A(_08966_),
    .B(_08970_),
    .X(_08971_));
 sky130_fd_sc_hd__and2b_1 _16392_ (.A_N(_08959_),
    .B(_08971_),
    .X(_08972_));
 sky130_fd_sc_hd__and2b_1 _16393_ (.A_N(_08971_),
    .B(_08959_),
    .X(_08973_));
 sky130_fd_sc_hd__nor2_1 _16394_ (.A(_08972_),
    .B(_08973_),
    .Y(_08974_));
 sky130_fd_sc_hd__clkbuf_4 _16395_ (.A(_08897_),
    .X(_08975_));
 sky130_fd_sc_hd__a21o_1 _16396_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[9] ),
    .A2(_08975_),
    .B1(_08896_),
    .X(_08976_));
 sky130_fd_sc_hd__a31o_1 _16397_ (.A1(_08679_),
    .A2(_08688_),
    .A3(_08928_),
    .B1(_08929_),
    .X(_08977_));
 sky130_fd_sc_hd__xnor2_1 _16398_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[10] ),
    .B(_08897_),
    .Y(_08978_));
 sky130_fd_sc_hd__xnor2_1 _16399_ (.A(_08977_),
    .B(_08978_),
    .Y(_08979_));
 sky130_fd_sc_hd__xor2_1 _16400_ (.A(_08976_),
    .B(_08979_),
    .X(_08980_));
 sky130_fd_sc_hd__xnor2_1 _16401_ (.A(_08974_),
    .B(_08980_),
    .Y(_08981_));
 sky130_fd_sc_hd__and2b_1 _16402_ (.A_N(_08936_),
    .B(_08934_),
    .X(_08982_));
 sky130_fd_sc_hd__a21oi_1 _16403_ (.A1(_08937_),
    .A2(_08943_),
    .B1(_08982_),
    .Y(_08983_));
 sky130_fd_sc_hd__xnor2_1 _16404_ (.A(_08981_),
    .B(_08983_),
    .Y(_08984_));
 sky130_fd_sc_hd__a21oi_1 _16405_ (.A1(_08938_),
    .A2(_08942_),
    .B1(_08940_),
    .Y(_08985_));
 sky130_fd_sc_hd__xnor2_1 _16406_ (.A(_08984_),
    .B(_08985_),
    .Y(_08986_));
 sky130_fd_sc_hd__or2_1 _16407_ (.A(_08944_),
    .B(_08946_),
    .X(_08987_));
 sky130_fd_sc_hd__o21a_1 _16408_ (.A1(_08947_),
    .A2(_08948_),
    .B1(_08987_),
    .X(_08988_));
 sky130_fd_sc_hd__xor2_1 _16409_ (.A(_08986_),
    .B(_08988_),
    .X(_08989_));
 sky130_fd_sc_hd__and2_1 _16410_ (.A(_08952_),
    .B(_08989_),
    .X(_08990_));
 sky130_fd_sc_hd__nor2_1 _16411_ (.A(_08952_),
    .B(_08989_),
    .Y(_08991_));
 sky130_fd_sc_hd__nor2_1 _16412_ (.A(_08990_),
    .B(_08991_),
    .Y(_08992_));
 sky130_fd_sc_hd__a21oi_1 _16413_ (.A1(_08920_),
    .A2(_08914_),
    .B1(_08954_),
    .Y(_08993_));
 sky130_fd_sc_hd__a31o_1 _16414_ (.A1(_08872_),
    .A2(_08916_),
    .A3(_08955_),
    .B1(_08993_),
    .X(_08994_));
 sky130_fd_sc_hd__nand2_1 _16415_ (.A(_08992_),
    .B(_08994_),
    .Y(_08995_));
 sky130_fd_sc_hd__o21a_1 _16416_ (.A1(_08992_),
    .A2(_08994_),
    .B1(_08265_),
    .X(_08996_));
 sky130_fd_sc_hd__a22o_1 _16417_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[10] ),
    .A2(_08066_),
    .B1(_08995_),
    .B2(_08996_),
    .X(_08997_));
 sky130_fd_sc_hd__and2_1 _16418_ (.A(_08831_),
    .B(_08997_),
    .X(_08998_));
 sky130_fd_sc_hd__clkbuf_1 _16419_ (.A(_08998_),
    .X(_00542_));
 sky130_fd_sc_hd__inv_2 _16420_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[11] ),
    .Y(_08999_));
 sky130_fd_sc_hd__nor2_1 _16421_ (.A(_08986_),
    .B(_08988_),
    .Y(_09000_));
 sky130_fd_sc_hd__nor2_1 _16422_ (.A(_08981_),
    .B(_08983_),
    .Y(_09001_));
 sky130_fd_sc_hd__nor2_1 _16423_ (.A(_08984_),
    .B(_08985_),
    .Y(_09002_));
 sky130_fd_sc_hd__or2b_1 _16424_ (.A(_08965_),
    .B_N(_08964_),
    .X(_09003_));
 sky130_fd_sc_hd__nand2_1 _16425_ (.A(_08966_),
    .B(_08970_),
    .Y(_09004_));
 sky130_fd_sc_hd__o21ai_1 _16426_ (.A1(_08693_),
    .A2(_08690_),
    .B1(_08679_),
    .Y(_09005_));
 sky130_fd_sc_hd__nor2_2 _16427_ (.A(_08967_),
    .B(_09005_),
    .Y(_09006_));
 sky130_fd_sc_hd__xnor2_4 _16428_ (.A(_08932_),
    .B(_09006_),
    .Y(_09007_));
 sky130_fd_sc_hd__and4b_1 _16429_ (.A_N(\top_inst.grid_inst.data_path_wires[8][4] ),
    .B(\top_inst.grid_inst.data_path_wires[8][5] ),
    .C(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[6] ),
    .D(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[7] ),
    .X(_09008_));
 sky130_fd_sc_hd__a2bb2o_1 _16430_ (.A1_N(_08876_),
    .A2_N(\top_inst.grid_inst.data_path_wires[8][4] ),
    .B1(\top_inst.grid_inst.data_path_wires[8][5] ),
    .B2(_08697_),
    .X(_09009_));
 sky130_fd_sc_hd__and2b_1 _16431_ (.A_N(_09008_),
    .B(_09009_),
    .X(_09010_));
 sky130_fd_sc_hd__nand2_1 _16432_ (.A(_08676_),
    .B(_08695_),
    .Y(_09011_));
 sky130_fd_sc_hd__xnor2_1 _16433_ (.A(_09010_),
    .B(_09011_),
    .Y(_09012_));
 sky130_fd_sc_hd__o21ba_1 _16434_ (.A1(_08961_),
    .A2(_08963_),
    .B1_N(_08960_),
    .X(_09013_));
 sky130_fd_sc_hd__xnor2_1 _16435_ (.A(_09012_),
    .B(_09013_),
    .Y(_09014_));
 sky130_fd_sc_hd__nand2_1 _16436_ (.A(_09007_),
    .B(_09014_),
    .Y(_09015_));
 sky130_fd_sc_hd__or2_1 _16437_ (.A(_09007_),
    .B(_09014_),
    .X(_09016_));
 sky130_fd_sc_hd__nand2_1 _16438_ (.A(_09015_),
    .B(_09016_),
    .Y(_09017_));
 sky130_fd_sc_hd__a21oi_1 _16439_ (.A1(_09003_),
    .A2(_09004_),
    .B1(_09017_),
    .Y(_09018_));
 sky130_fd_sc_hd__nand3_1 _16440_ (.A(_09003_),
    .B(_09004_),
    .C(_09017_),
    .Y(_09019_));
 sky130_fd_sc_hd__or2b_1 _16441_ (.A(_09018_),
    .B_N(_09019_),
    .X(_09020_));
 sky130_fd_sc_hd__a21o_1 _16442_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[10] ),
    .A2(_08975_),
    .B1(_08896_),
    .X(_09021_));
 sky130_fd_sc_hd__a32o_1 _16443_ (.A1(_08679_),
    .A2(_08688_),
    .A3(_08968_),
    .B1(_08967_),
    .B2(_08677_),
    .X(_09022_));
 sky130_fd_sc_hd__xnor2_1 _16444_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[11] ),
    .B(_08897_),
    .Y(_09023_));
 sky130_fd_sc_hd__xnor2_1 _16445_ (.A(_09022_),
    .B(_09023_),
    .Y(_09024_));
 sky130_fd_sc_hd__xor2_1 _16446_ (.A(_09021_),
    .B(_09024_),
    .X(_09025_));
 sky130_fd_sc_hd__xnor2_1 _16447_ (.A(_09020_),
    .B(_09025_),
    .Y(_09026_));
 sky130_fd_sc_hd__a21o_1 _16448_ (.A1(_08974_),
    .A2(_08980_),
    .B1(_08972_),
    .X(_09027_));
 sky130_fd_sc_hd__xnor2_1 _16449_ (.A(_09026_),
    .B(_09027_),
    .Y(_09028_));
 sky130_fd_sc_hd__or2b_1 _16450_ (.A(_08978_),
    .B_N(_08977_),
    .X(_09029_));
 sky130_fd_sc_hd__a21bo_1 _16451_ (.A1(_08976_),
    .A2(_08979_),
    .B1_N(_09029_),
    .X(_09030_));
 sky130_fd_sc_hd__xnor2_1 _16452_ (.A(_09028_),
    .B(_09030_),
    .Y(_09031_));
 sky130_fd_sc_hd__o21ai_2 _16453_ (.A1(_09001_),
    .A2(_09002_),
    .B1(_09031_),
    .Y(_09032_));
 sky130_fd_sc_hd__or3_1 _16454_ (.A(_09001_),
    .B(_09002_),
    .C(_09031_),
    .X(_09033_));
 sky130_fd_sc_hd__and2_1 _16455_ (.A(_09032_),
    .B(_09033_),
    .X(_09034_));
 sky130_fd_sc_hd__xnor2_1 _16456_ (.A(_09000_),
    .B(_09034_),
    .Y(_09035_));
 sky130_fd_sc_hd__a21oi_1 _16457_ (.A1(_08992_),
    .A2(_08994_),
    .B1(_08990_),
    .Y(_09036_));
 sky130_fd_sc_hd__xnor2_1 _16458_ (.A(_09035_),
    .B(_09036_),
    .Y(_09037_));
 sky130_fd_sc_hd__mux2_1 _16459_ (.A0(_08999_),
    .A1(_09037_),
    .S(_05335_),
    .X(_09038_));
 sky130_fd_sc_hd__nor2_1 _16460_ (.A(_05440_),
    .B(_09038_),
    .Y(_00543_));
 sky130_fd_sc_hd__or2b_1 _16461_ (.A(_09013_),
    .B_N(_09012_),
    .X(_09039_));
 sky130_fd_sc_hd__nand2_2 _16462_ (.A(_08679_),
    .B(_08695_),
    .Y(_09040_));
 sky130_fd_sc_hd__nor2_1 _16463_ (.A(_08876_),
    .B(_08673_),
    .Y(_09041_));
 sky130_fd_sc_hd__and3_1 _16464_ (.A(_08697_),
    .B(_08676_),
    .C(_09041_),
    .X(_09042_));
 sky130_fd_sc_hd__a21oi_1 _16465_ (.A1(_08697_),
    .A2(_08676_),
    .B1(_09041_),
    .Y(_09043_));
 sky130_fd_sc_hd__or2_1 _16466_ (.A(_09042_),
    .B(_09043_),
    .X(_09044_));
 sky130_fd_sc_hd__xor2_1 _16467_ (.A(_09040_),
    .B(_09044_),
    .X(_09045_));
 sky130_fd_sc_hd__a31o_1 _16468_ (.A1(_08677_),
    .A2(_08695_),
    .A3(_09009_),
    .B1(_09008_),
    .X(_09046_));
 sky130_fd_sc_hd__xor2_1 _16469_ (.A(_09045_),
    .B(_09046_),
    .X(_09047_));
 sky130_fd_sc_hd__nand2_1 _16470_ (.A(_09007_),
    .B(_09047_),
    .Y(_09048_));
 sky130_fd_sc_hd__or2_1 _16471_ (.A(_09007_),
    .B(_09047_),
    .X(_09049_));
 sky130_fd_sc_hd__nand2_1 _16472_ (.A(_09048_),
    .B(_09049_),
    .Y(_09050_));
 sky130_fd_sc_hd__a21o_1 _16473_ (.A1(_09039_),
    .A2(_09015_),
    .B1(_09050_),
    .X(_09051_));
 sky130_fd_sc_hd__nand3_1 _16474_ (.A(_09039_),
    .B(_09015_),
    .C(_09050_),
    .Y(_09052_));
 sky130_fd_sc_hd__nand2_1 _16475_ (.A(_09051_),
    .B(_09052_),
    .Y(_09053_));
 sky130_fd_sc_hd__a21o_1 _16476_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[11] ),
    .A2(_08975_),
    .B1(_08896_),
    .X(_09054_));
 sky130_fd_sc_hd__o21ba_2 _16477_ (.A1(_08932_),
    .A2(_09005_),
    .B1_N(_08967_),
    .X(_09055_));
 sky130_fd_sc_hd__xnor2_1 _16478_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[12] ),
    .B(_08897_),
    .Y(_09056_));
 sky130_fd_sc_hd__nor2_1 _16479_ (.A(_09055_),
    .B(_09056_),
    .Y(_09057_));
 sky130_fd_sc_hd__and2_1 _16480_ (.A(_09055_),
    .B(_09056_),
    .X(_09058_));
 sky130_fd_sc_hd__nor2_1 _16481_ (.A(_09057_),
    .B(_09058_),
    .Y(_09059_));
 sky130_fd_sc_hd__xnor2_2 _16482_ (.A(_09054_),
    .B(_09059_),
    .Y(_09060_));
 sky130_fd_sc_hd__xor2_1 _16483_ (.A(_09053_),
    .B(_09060_),
    .X(_09061_));
 sky130_fd_sc_hd__a21o_1 _16484_ (.A1(_09019_),
    .A2(_09025_),
    .B1(_09018_),
    .X(_09062_));
 sky130_fd_sc_hd__xnor2_1 _16485_ (.A(_09061_),
    .B(_09062_),
    .Y(_09063_));
 sky130_fd_sc_hd__or2b_1 _16486_ (.A(_09023_),
    .B_N(_09022_),
    .X(_09064_));
 sky130_fd_sc_hd__a21bo_1 _16487_ (.A1(_09021_),
    .A2(_09024_),
    .B1_N(_09064_),
    .X(_09065_));
 sky130_fd_sc_hd__xnor2_1 _16488_ (.A(_09063_),
    .B(_09065_),
    .Y(_09066_));
 sky130_fd_sc_hd__or2b_1 _16489_ (.A(_09028_),
    .B_N(_09030_),
    .X(_09067_));
 sky130_fd_sc_hd__a21bo_1 _16490_ (.A1(_09026_),
    .A2(_09027_),
    .B1_N(_09067_),
    .X(_09068_));
 sky130_fd_sc_hd__and2_1 _16491_ (.A(_09066_),
    .B(_09068_),
    .X(_09069_));
 sky130_fd_sc_hd__nor2_1 _16492_ (.A(_09066_),
    .B(_09068_),
    .Y(_09070_));
 sky130_fd_sc_hd__nor2_1 _16493_ (.A(_09069_),
    .B(_09070_),
    .Y(_09071_));
 sky130_fd_sc_hd__xor2_2 _16494_ (.A(_09032_),
    .B(_09071_),
    .X(_09072_));
 sky130_fd_sc_hd__nand2_1 _16495_ (.A(_09000_),
    .B(_09034_),
    .Y(_09073_));
 sky130_fd_sc_hd__o21a_1 _16496_ (.A1(_09035_),
    .A2(_09036_),
    .B1(_09073_),
    .X(_09074_));
 sky130_fd_sc_hd__nor2_1 _16497_ (.A(_09072_),
    .B(_09074_),
    .Y(_09075_));
 sky130_fd_sc_hd__a21o_1 _16498_ (.A1(_09072_),
    .A2(_09074_),
    .B1(_05353_),
    .X(_09076_));
 sky130_fd_sc_hd__a2bb2o_1 _16499_ (.A1_N(_09075_),
    .A2_N(_09076_),
    .B1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[12] ),
    .B2(_07816_),
    .X(_09077_));
 sky130_fd_sc_hd__and2_1 _16500_ (.A(_08831_),
    .B(_09077_),
    .X(_09078_));
 sky130_fd_sc_hd__clkbuf_1 _16501_ (.A(_09078_),
    .X(_00544_));
 sky130_fd_sc_hd__nand2_1 _16502_ (.A(net1008),
    .B(_05403_),
    .Y(_09079_));
 sky130_fd_sc_hd__nand2_1 _16503_ (.A(_09045_),
    .B(_09046_),
    .Y(_09080_));
 sky130_fd_sc_hd__nand2_1 _16504_ (.A(_08679_),
    .B(_08697_),
    .Y(_09081_));
 sky130_fd_sc_hd__o21a_1 _16505_ (.A1(_08876_),
    .A2(_08677_),
    .B1(_09081_),
    .X(_09082_));
 sky130_fd_sc_hd__nor3_1 _16506_ (.A(_08876_),
    .B(_08677_),
    .C(_09081_),
    .Y(_09083_));
 sky130_fd_sc_hd__nor2_1 _16507_ (.A(_09082_),
    .B(_09083_),
    .Y(_09084_));
 sky130_fd_sc_hd__xnor2_1 _16508_ (.A(_09040_),
    .B(_09084_),
    .Y(_09085_));
 sky130_fd_sc_hd__o21ba_1 _16509_ (.A1(_09040_),
    .A2(_09043_),
    .B1_N(_09042_),
    .X(_09086_));
 sky130_fd_sc_hd__xnor2_1 _16510_ (.A(_09085_),
    .B(_09086_),
    .Y(_09087_));
 sky130_fd_sc_hd__nand2_1 _16511_ (.A(_09007_),
    .B(_09087_),
    .Y(_09088_));
 sky130_fd_sc_hd__or2_1 _16512_ (.A(_09007_),
    .B(_09087_),
    .X(_09089_));
 sky130_fd_sc_hd__nand2_1 _16513_ (.A(_09088_),
    .B(_09089_),
    .Y(_09090_));
 sky130_fd_sc_hd__a21o_1 _16514_ (.A1(_09080_),
    .A2(_09048_),
    .B1(_09090_),
    .X(_09091_));
 sky130_fd_sc_hd__nand3_1 _16515_ (.A(_09080_),
    .B(_09048_),
    .C(_09090_),
    .Y(_09092_));
 sky130_fd_sc_hd__a21o_1 _16516_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[12] ),
    .A2(_08975_),
    .B1(_08896_),
    .X(_09093_));
 sky130_fd_sc_hd__xnor2_1 _16517_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[13] ),
    .B(_08975_),
    .Y(_09094_));
 sky130_fd_sc_hd__nor2_1 _16518_ (.A(_09055_),
    .B(_09094_),
    .Y(_09095_));
 sky130_fd_sc_hd__and2_1 _16519_ (.A(_09055_),
    .B(_09094_),
    .X(_09096_));
 sky130_fd_sc_hd__nor2_1 _16520_ (.A(_09095_),
    .B(_09096_),
    .Y(_09097_));
 sky130_fd_sc_hd__xor2_1 _16521_ (.A(_09093_),
    .B(_09097_),
    .X(_09098_));
 sky130_fd_sc_hd__and3_1 _16522_ (.A(_09091_),
    .B(_09092_),
    .C(_09098_),
    .X(_09099_));
 sky130_fd_sc_hd__a21oi_1 _16523_ (.A1(_09091_),
    .A2(_09092_),
    .B1(_09098_),
    .Y(_09100_));
 sky130_fd_sc_hd__nor2_1 _16524_ (.A(_09099_),
    .B(_09100_),
    .Y(_09101_));
 sky130_fd_sc_hd__o21ai_2 _16525_ (.A1(_09053_),
    .A2(_09060_),
    .B1(_09051_),
    .Y(_09102_));
 sky130_fd_sc_hd__xnor2_1 _16526_ (.A(_09101_),
    .B(_09102_),
    .Y(_09103_));
 sky130_fd_sc_hd__a21o_1 _16527_ (.A1(_09054_),
    .A2(_09059_),
    .B1(_09057_),
    .X(_09104_));
 sky130_fd_sc_hd__xnor2_1 _16528_ (.A(_09103_),
    .B(_09104_),
    .Y(_09105_));
 sky130_fd_sc_hd__or2b_1 _16529_ (.A(_09063_),
    .B_N(_09065_),
    .X(_09106_));
 sky130_fd_sc_hd__a21bo_1 _16530_ (.A1(_09061_),
    .A2(_09062_),
    .B1_N(_09106_),
    .X(_09107_));
 sky130_fd_sc_hd__nand2_1 _16531_ (.A(_09105_),
    .B(_09107_),
    .Y(_09108_));
 sky130_fd_sc_hd__or2_1 _16532_ (.A(_09105_),
    .B(_09107_),
    .X(_09109_));
 sky130_fd_sc_hd__and2_1 _16533_ (.A(_09108_),
    .B(_09109_),
    .X(_09110_));
 sky130_fd_sc_hd__xor2_1 _16534_ (.A(_09069_),
    .B(_09110_),
    .X(_09111_));
 sky130_fd_sc_hd__and2b_1 _16535_ (.A_N(_09032_),
    .B(_09071_),
    .X(_09112_));
 sky130_fd_sc_hd__o21bai_2 _16536_ (.A1(_09072_),
    .A2(_09074_),
    .B1_N(_09112_),
    .Y(_09113_));
 sky130_fd_sc_hd__a21oi_1 _16537_ (.A1(_09111_),
    .A2(_09113_),
    .B1(_05406_),
    .Y(_09114_));
 sky130_fd_sc_hd__o21ai_1 _16538_ (.A1(_09111_),
    .A2(_09113_),
    .B1(_09114_),
    .Y(_09115_));
 sky130_fd_sc_hd__a21oi_1 _16539_ (.A1(_09079_),
    .A2(_09115_),
    .B1(_04867_),
    .Y(_00545_));
 sky130_fd_sc_hd__a21oi_1 _16540_ (.A1(_09080_),
    .A2(_09048_),
    .B1(_09090_),
    .Y(_09116_));
 sky130_fd_sc_hd__or2b_1 _16541_ (.A(_09086_),
    .B_N(_09085_),
    .X(_09117_));
 sky130_fd_sc_hd__and3_1 _16542_ (.A(_08679_),
    .B(_08697_),
    .C(_08695_),
    .X(_09118_));
 sky130_fd_sc_hd__o21ba_1 _16543_ (.A1(_09040_),
    .A2(_09082_),
    .B1_N(_09083_),
    .X(_09119_));
 sky130_fd_sc_hd__o21a_1 _16544_ (.A1(_08876_),
    .A2(_08679_),
    .B1(_09081_),
    .X(_09120_));
 sky130_fd_sc_hd__a2bb2o_1 _16545_ (.A1_N(_09118_),
    .A2_N(_09119_),
    .B1(_09040_),
    .B2(_09120_),
    .X(_09121_));
 sky130_fd_sc_hd__xor2_1 _16546_ (.A(_09007_),
    .B(_09121_),
    .X(_09122_));
 sky130_fd_sc_hd__a21oi_1 _16547_ (.A1(_09117_),
    .A2(_09088_),
    .B1(_09122_),
    .Y(_09123_));
 sky130_fd_sc_hd__nand3_1 _16548_ (.A(_09117_),
    .B(_09088_),
    .C(_09122_),
    .Y(_09124_));
 sky130_fd_sc_hd__or2b_1 _16549_ (.A(_09123_),
    .B_N(_09124_),
    .X(_09125_));
 sky130_fd_sc_hd__a21oi_1 _16550_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[13] ),
    .A2(_08975_),
    .B1(_08896_),
    .Y(_09126_));
 sky130_fd_sc_hd__xnor2_1 _16551_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[14] ),
    .B(_08975_),
    .Y(_09127_));
 sky130_fd_sc_hd__nor2_1 _16552_ (.A(_09055_),
    .B(_09127_),
    .Y(_09128_));
 sky130_fd_sc_hd__and2_1 _16553_ (.A(_09055_),
    .B(_09127_),
    .X(_09129_));
 sky130_fd_sc_hd__nor2_1 _16554_ (.A(_09128_),
    .B(_09129_),
    .Y(_09130_));
 sky130_fd_sc_hd__xnor2_1 _16555_ (.A(_09126_),
    .B(_09130_),
    .Y(_09131_));
 sky130_fd_sc_hd__xnor2_1 _16556_ (.A(_09125_),
    .B(_09131_),
    .Y(_09132_));
 sky130_fd_sc_hd__o21ai_1 _16557_ (.A1(_09116_),
    .A2(_09099_),
    .B1(_09132_),
    .Y(_09133_));
 sky130_fd_sc_hd__or3_1 _16558_ (.A(_09116_),
    .B(_09099_),
    .C(_09132_),
    .X(_09134_));
 sky130_fd_sc_hd__nand2_1 _16559_ (.A(_09133_),
    .B(_09134_),
    .Y(_09135_));
 sky130_fd_sc_hd__a21oi_2 _16560_ (.A1(_09093_),
    .A2(_09097_),
    .B1(_09095_),
    .Y(_09136_));
 sky130_fd_sc_hd__xnor2_2 _16561_ (.A(_09135_),
    .B(_09136_),
    .Y(_09137_));
 sky130_fd_sc_hd__or2b_1 _16562_ (.A(_09103_),
    .B_N(_09104_),
    .X(_09138_));
 sky130_fd_sc_hd__a21boi_2 _16563_ (.A1(_09101_),
    .A2(_09102_),
    .B1_N(_09138_),
    .Y(_09139_));
 sky130_fd_sc_hd__xnor2_1 _16564_ (.A(_09137_),
    .B(_09139_),
    .Y(_09140_));
 sky130_fd_sc_hd__nor2_1 _16565_ (.A(_09108_),
    .B(_09140_),
    .Y(_09141_));
 sky130_fd_sc_hd__and2_1 _16566_ (.A(_09108_),
    .B(_09140_),
    .X(_09142_));
 sky130_fd_sc_hd__nor2_1 _16567_ (.A(_09141_),
    .B(_09142_),
    .Y(_09143_));
 sky130_fd_sc_hd__a32o_1 _16568_ (.A1(_09066_),
    .A2(_09068_),
    .A3(_09110_),
    .B1(_09111_),
    .B2(_09113_),
    .X(_09144_));
 sky130_fd_sc_hd__nand2_1 _16569_ (.A(_09143_),
    .B(_09144_),
    .Y(_09145_));
 sky130_fd_sc_hd__o21a_1 _16570_ (.A1(_09143_),
    .A2(_09144_),
    .B1(_08265_),
    .X(_09146_));
 sky130_fd_sc_hd__a22o_1 _16571_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[14] ),
    .A2(_08066_),
    .B1(_09145_),
    .B2(_09146_),
    .X(_09147_));
 sky130_fd_sc_hd__and2_1 _16572_ (.A(_08831_),
    .B(_09147_),
    .X(_09148_));
 sky130_fd_sc_hd__clkbuf_1 _16573_ (.A(_09148_),
    .X(_00546_));
 sky130_fd_sc_hd__and2_1 _16574_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[15] ),
    .B(_05634_),
    .X(_09149_));
 sky130_fd_sc_hd__a21oi_1 _16575_ (.A1(_09124_),
    .A2(_09131_),
    .B1(_09123_),
    .Y(_09150_));
 sky130_fd_sc_hd__and2b_1 _16576_ (.A_N(_09007_),
    .B(_09121_),
    .X(_09151_));
 sky130_fd_sc_hd__a21o_1 _16577_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[14] ),
    .A2(_08975_),
    .B1(_08896_),
    .X(_09152_));
 sky130_fd_sc_hd__xnor2_2 _16578_ (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[15] ),
    .B(_08975_),
    .Y(_09153_));
 sky130_fd_sc_hd__xnor2_1 _16579_ (.A(_09055_),
    .B(_09153_),
    .Y(_09154_));
 sky130_fd_sc_hd__xnor2_1 _16580_ (.A(_09152_),
    .B(_09154_),
    .Y(_09155_));
 sky130_fd_sc_hd__or2_1 _16581_ (.A(_09151_),
    .B(_09155_),
    .X(_09156_));
 sky130_fd_sc_hd__nand2_1 _16582_ (.A(_09151_),
    .B(_09155_),
    .Y(_09157_));
 sky130_fd_sc_hd__and2_1 _16583_ (.A(_09156_),
    .B(_09157_),
    .X(_09158_));
 sky130_fd_sc_hd__xnor2_1 _16584_ (.A(_09150_),
    .B(_09158_),
    .Y(_09159_));
 sky130_fd_sc_hd__o21ba_1 _16585_ (.A1(_09126_),
    .A2(_09129_),
    .B1_N(_09128_),
    .X(_09160_));
 sky130_fd_sc_hd__xnor2_1 _16586_ (.A(_09159_),
    .B(_09160_),
    .Y(_09161_));
 sky130_fd_sc_hd__o21a_1 _16587_ (.A1(_09135_),
    .A2(_09136_),
    .B1(_09133_),
    .X(_09162_));
 sky130_fd_sc_hd__or2_1 _16588_ (.A(_09161_),
    .B(_09162_),
    .X(_09163_));
 sky130_fd_sc_hd__nand2_1 _16589_ (.A(_09161_),
    .B(_09162_),
    .Y(_09164_));
 sky130_fd_sc_hd__and4bb_1 _16590_ (.A_N(_09137_),
    .B_N(_09139_),
    .C(_09163_),
    .D(_09164_),
    .X(_09165_));
 sky130_fd_sc_hd__and2_1 _16591_ (.A(_09163_),
    .B(_09164_),
    .X(_09166_));
 sky130_fd_sc_hd__o21ba_1 _16592_ (.A1(_09137_),
    .A2(_09139_),
    .B1_N(_09166_),
    .X(_09167_));
 sky130_fd_sc_hd__a21oi_1 _16593_ (.A1(_09143_),
    .A2(_09144_),
    .B1(_09141_),
    .Y(_09168_));
 sky130_fd_sc_hd__nor2_1 _16594_ (.A(_09165_),
    .B(_09167_),
    .Y(_09169_));
 sky130_fd_sc_hd__a211o_1 _16595_ (.A1(_09143_),
    .A2(_09144_),
    .B1(_09169_),
    .C1(_09141_),
    .X(_09170_));
 sky130_fd_sc_hd__o311a_1 _16596_ (.A1(_09165_),
    .A2(_09167_),
    .A3(_09168_),
    .B1(_09170_),
    .C1(_05313_),
    .X(_09171_));
 sky130_fd_sc_hd__o21a_1 _16597_ (.A1(_09149_),
    .A2(_09171_),
    .B1(_04870_),
    .X(_00547_));
 sky130_fd_sc_hd__or2_1 _16598_ (.A(_09150_),
    .B(_09158_),
    .X(_09172_));
 sky130_fd_sc_hd__o21a_1 _16599_ (.A1(_09159_),
    .A2(_09160_),
    .B1(_09172_),
    .X(_09173_));
 sky130_fd_sc_hd__xnor2_1 _16600_ (.A(_09156_),
    .B(_09173_),
    .Y(_09174_));
 sky130_fd_sc_hd__a21o_1 _16601_ (.A1(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[15] ),
    .A2(_08975_),
    .B1(_08896_),
    .X(_09175_));
 sky130_fd_sc_hd__o21a_1 _16602_ (.A1(_09055_),
    .A2(_09153_),
    .B1(_09152_),
    .X(_09176_));
 sky130_fd_sc_hd__a21oi_1 _16603_ (.A1(_09055_),
    .A2(_09153_),
    .B1(_09176_),
    .Y(_09177_));
 sky130_fd_sc_hd__xnor2_1 _16604_ (.A(_09163_),
    .B(_09177_),
    .Y(_09178_));
 sky130_fd_sc_hd__xnor2_1 _16605_ (.A(_09175_),
    .B(_09178_),
    .Y(_09179_));
 sky130_fd_sc_hd__xnor2_1 _16606_ (.A(_09174_),
    .B(_09179_),
    .Y(_09180_));
 sky130_fd_sc_hd__nor2_1 _16607_ (.A(_09165_),
    .B(_09180_),
    .Y(_09181_));
 sky130_fd_sc_hd__o31a_1 _16608_ (.A1(_09165_),
    .A2(_09167_),
    .A3(_09168_),
    .B1(_09181_),
    .X(_09182_));
 sky130_fd_sc_hd__or2_1 _16609_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[16] ),
    .B(_07866_),
    .X(_09183_));
 sky130_fd_sc_hd__clkbuf_4 _16610_ (.A(_07617_),
    .X(_09184_));
 sky130_fd_sc_hd__o211a_1 _16611_ (.A1(_08870_),
    .A2(_09182_),
    .B1(_09183_),
    .C1(_09184_),
    .X(_00548_));
 sky130_fd_sc_hd__clkbuf_4 _16612_ (.A(_05269_),
    .X(_09185_));
 sky130_fd_sc_hd__mux2_4 _16613_ (.A0(\top_inst.skew_buff_inst.row[2].output_reg[0] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[16] ),
    .S(_07059_),
    .X(_09186_));
 sky130_fd_sc_hd__buf_2 _16614_ (.A(_09186_),
    .X(_09187_));
 sky130_fd_sc_hd__clkbuf_4 _16615_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[0] ),
    .X(_09188_));
 sky130_fd_sc_hd__clkbuf_4 _16616_ (.A(_09188_),
    .X(_09189_));
 sky130_fd_sc_hd__or2_1 _16617_ (.A(_09189_),
    .B(_08684_),
    .X(_09190_));
 sky130_fd_sc_hd__o211a_1 _16618_ (.A1(_09185_),
    .A2(_09187_),
    .B1(_09190_),
    .C1(_09184_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_4 _16619_ (.A0(\top_inst.skew_buff_inst.row[2].output_reg[1] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[17] ),
    .S(_07059_),
    .X(_09191_));
 sky130_fd_sc_hd__clkbuf_4 _16620_ (.A(net1119),
    .X(_09192_));
 sky130_fd_sc_hd__clkbuf_4 _16621_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[1] ),
    .X(_09193_));
 sky130_fd_sc_hd__clkbuf_4 _16622_ (.A(_09193_),
    .X(_09194_));
 sky130_fd_sc_hd__or2_1 _16623_ (.A(_09194_),
    .B(_08684_),
    .X(_09195_));
 sky130_fd_sc_hd__o211a_1 _16624_ (.A1(_09185_),
    .A2(_09192_),
    .B1(_09195_),
    .C1(_09184_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_4 _16625_ (.A0(\top_inst.skew_buff_inst.row[2].output_reg[2] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[18] ),
    .S(_07059_),
    .X(_09196_));
 sky130_fd_sc_hd__clkbuf_4 _16626_ (.A(net224),
    .X(_09197_));
 sky130_fd_sc_hd__clkbuf_4 _16627_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[2] ),
    .X(_09198_));
 sky130_fd_sc_hd__clkbuf_4 _16628_ (.A(_05772_),
    .X(_09199_));
 sky130_fd_sc_hd__or2_1 _16629_ (.A(_09198_),
    .B(_09199_),
    .X(_09200_));
 sky130_fd_sc_hd__o211a_1 _16630_ (.A1(_09185_),
    .A2(_09197_),
    .B1(_09200_),
    .C1(_09184_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_4 _16631_ (.A0(\top_inst.skew_buff_inst.row[2].output_reg[3] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[19] ),
    .S(_07059_),
    .X(_09201_));
 sky130_fd_sc_hd__clkbuf_4 _16632_ (.A(_09201_),
    .X(_09202_));
 sky130_fd_sc_hd__buf_4 _16633_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[3] ),
    .X(_09203_));
 sky130_fd_sc_hd__or2_1 _16634_ (.A(_09203_),
    .B(_09199_),
    .X(_09204_));
 sky130_fd_sc_hd__o211a_1 _16635_ (.A1(_09185_),
    .A2(_09202_),
    .B1(_09204_),
    .C1(_09184_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_4 _16636_ (.A0(\top_inst.skew_buff_inst.row[2].output_reg[4] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[20] ),
    .S(_05265_),
    .X(_09205_));
 sky130_fd_sc_hd__buf_4 _16637_ (.A(net216),
    .X(_09206_));
 sky130_fd_sc_hd__clkbuf_4 _16638_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[4] ),
    .X(_09207_));
 sky130_fd_sc_hd__or2_1 _16639_ (.A(_09207_),
    .B(_09199_),
    .X(_09208_));
 sky130_fd_sc_hd__o211a_1 _16640_ (.A1(_09185_),
    .A2(_09206_),
    .B1(_09208_),
    .C1(_09184_),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_4 _16641_ (.A0(\top_inst.skew_buff_inst.row[2].output_reg[5] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[21] ),
    .S(_05265_),
    .X(_09209_));
 sky130_fd_sc_hd__clkbuf_4 _16642_ (.A(_09209_),
    .X(_09210_));
 sky130_fd_sc_hd__buf_2 _16643_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[5] ),
    .X(_09211_));
 sky130_fd_sc_hd__or2_1 _16644_ (.A(_09211_),
    .B(_09199_),
    .X(_09212_));
 sky130_fd_sc_hd__o211a_1 _16645_ (.A1(_09185_),
    .A2(_09210_),
    .B1(_09212_),
    .C1(_09184_),
    .X(_00554_));
 sky130_fd_sc_hd__buf_2 _16646_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[6] ),
    .X(_09213_));
 sky130_fd_sc_hd__mux2_4 _16647_ (.A0(\top_inst.skew_buff_inst.row[2].output_reg[6] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[22] ),
    .S(_05266_),
    .X(_09214_));
 sky130_fd_sc_hd__buf_2 _16648_ (.A(_09214_),
    .X(_09215_));
 sky130_fd_sc_hd__or2_1 _16649_ (.A(_05269_),
    .B(_09215_),
    .X(_09216_));
 sky130_fd_sc_hd__o211a_1 _16650_ (.A1(_09213_),
    .A2(_05276_),
    .B1(_09216_),
    .C1(_09184_),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_2 _16651_ (.A0(\top_inst.skew_buff_inst.row[2].output_reg[7] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[23] ),
    .S(net185),
    .X(_09217_));
 sky130_fd_sc_hd__buf_6 _16652_ (.A(_09217_),
    .X(_09218_));
 sky130_fd_sc_hd__clkbuf_4 _16653_ (.A(net219),
    .X(_09219_));
 sky130_fd_sc_hd__or2_1 _16654_ (.A(_05269_),
    .B(_09219_),
    .X(_09220_));
 sky130_fd_sc_hd__o211a_1 _16655_ (.A1(net1058),
    .A2(_05276_),
    .B1(_09220_),
    .C1(_09184_),
    .X(_00556_));
 sky130_fd_sc_hd__a21oi_1 _16656_ (.A1(_09189_),
    .A2(_09187_),
    .B1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[0] ),
    .Y(_09221_));
 sky130_fd_sc_hd__and3_1 _16657_ (.A(_09189_),
    .B(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[0] ),
    .C(_09187_),
    .X(_09222_));
 sky130_fd_sc_hd__o21ai_1 _16658_ (.A1(_09221_),
    .A2(_09222_),
    .B1(_08181_),
    .Y(_09223_));
 sky130_fd_sc_hd__o211a_1 _16659_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[0] ),
    .A2(_08183_),
    .B1(_09223_),
    .C1(_09184_),
    .X(_00557_));
 sky130_fd_sc_hd__a22o_1 _16660_ (.A1(_09194_),
    .A2(_09187_),
    .B1(_09192_),
    .B2(_09189_),
    .X(_09224_));
 sky130_fd_sc_hd__nand4_1 _16661_ (.A(_09194_),
    .B(_09189_),
    .C(_09187_),
    .D(_09192_),
    .Y(_09225_));
 sky130_fd_sc_hd__and3_1 _16662_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[1] ),
    .B(_09224_),
    .C(_09225_),
    .X(_09226_));
 sky130_fd_sc_hd__a21oi_1 _16663_ (.A1(_09224_),
    .A2(_09225_),
    .B1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[1] ),
    .Y(_09227_));
 sky130_fd_sc_hd__o21ba_1 _16664_ (.A1(_09226_),
    .A2(_09227_),
    .B1_N(_09222_),
    .X(_09228_));
 sky130_fd_sc_hd__nor3b_1 _16665_ (.A(_09226_),
    .B(_09227_),
    .C_N(_09222_),
    .Y(_09229_));
 sky130_fd_sc_hd__o21ai_1 _16666_ (.A1(_09228_),
    .A2(_09229_),
    .B1(_08181_),
    .Y(_09230_));
 sky130_fd_sc_hd__clkbuf_4 _16667_ (.A(_07617_),
    .X(_09231_));
 sky130_fd_sc_hd__o211a_1 _16668_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[1] ),
    .A2(_08183_),
    .B1(_09230_),
    .C1(_09231_),
    .X(_00558_));
 sky130_fd_sc_hd__nand2_1 _16669_ (.A(_09198_),
    .B(_09187_),
    .Y(_09232_));
 sky130_fd_sc_hd__a22o_1 _16670_ (.A1(_09194_),
    .A2(_09192_),
    .B1(_09197_),
    .B2(_09189_),
    .X(_09233_));
 sky130_fd_sc_hd__nand4_2 _16671_ (.A(_09194_),
    .B(_09189_),
    .C(_09192_),
    .D(_09197_),
    .Y(_09234_));
 sky130_fd_sc_hd__nand3_1 _16672_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[2] ),
    .B(_09233_),
    .C(_09234_),
    .Y(_09235_));
 sky130_fd_sc_hd__a21o_1 _16673_ (.A1(_09233_),
    .A2(_09234_),
    .B1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[2] ),
    .X(_09236_));
 sky130_fd_sc_hd__nand2_1 _16674_ (.A(_09235_),
    .B(_09236_),
    .Y(_09237_));
 sky130_fd_sc_hd__a21boi_1 _16675_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[1] ),
    .A2(_09224_),
    .B1_N(_09225_),
    .Y(_09238_));
 sky130_fd_sc_hd__xnor2_1 _16676_ (.A(_09237_),
    .B(_09238_),
    .Y(_09239_));
 sky130_fd_sc_hd__nor2_1 _16677_ (.A(_09232_),
    .B(_09239_),
    .Y(_09240_));
 sky130_fd_sc_hd__and2_1 _16678_ (.A(_09232_),
    .B(_09239_),
    .X(_09241_));
 sky130_fd_sc_hd__nor2_1 _16679_ (.A(_09240_),
    .B(_09241_),
    .Y(_09242_));
 sky130_fd_sc_hd__nand2_1 _16680_ (.A(_09229_),
    .B(_09242_),
    .Y(_09243_));
 sky130_fd_sc_hd__o21a_1 _16681_ (.A1(_09229_),
    .A2(_09242_),
    .B1(_08265_),
    .X(_09244_));
 sky130_fd_sc_hd__a22o_1 _16682_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[2] ),
    .A2(_08066_),
    .B1(_09243_),
    .B2(_09244_),
    .X(_09245_));
 sky130_fd_sc_hd__and2_1 _16683_ (.A(_08831_),
    .B(_09245_),
    .X(_09246_));
 sky130_fd_sc_hd__clkbuf_1 _16684_ (.A(_09246_),
    .X(_00559_));
 sky130_fd_sc_hd__nor2_1 _16685_ (.A(_09237_),
    .B(_09238_),
    .Y(_09247_));
 sky130_fd_sc_hd__a22o_1 _16686_ (.A1(_09194_),
    .A2(_09197_),
    .B1(_09202_),
    .B2(_09188_),
    .X(_09248_));
 sky130_fd_sc_hd__nand4_1 _16687_ (.A(_09194_),
    .B(_09188_),
    .C(_09197_),
    .D(_09202_),
    .Y(_09249_));
 sky130_fd_sc_hd__nand2_1 _16688_ (.A(_09248_),
    .B(_09249_),
    .Y(_09250_));
 sky130_fd_sc_hd__xnor2_1 _16689_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[3] ),
    .B(_09250_),
    .Y(_09251_));
 sky130_fd_sc_hd__nand2_1 _16690_ (.A(_09234_),
    .B(_09235_),
    .Y(_09252_));
 sky130_fd_sc_hd__xnor2_1 _16691_ (.A(_09251_),
    .B(_09252_),
    .Y(_09253_));
 sky130_fd_sc_hd__a22o_1 _16692_ (.A1(_09203_),
    .A2(_09187_),
    .B1(_09192_),
    .B2(_09198_),
    .X(_09254_));
 sky130_fd_sc_hd__nand4_2 _16693_ (.A(_09203_),
    .B(_09198_),
    .C(_09186_),
    .D(_09192_),
    .Y(_09255_));
 sky130_fd_sc_hd__and2_1 _16694_ (.A(_09254_),
    .B(_09255_),
    .X(_09256_));
 sky130_fd_sc_hd__xnor2_1 _16695_ (.A(_09253_),
    .B(_09256_),
    .Y(_09257_));
 sky130_fd_sc_hd__o21a_1 _16696_ (.A1(_09247_),
    .A2(_09240_),
    .B1(_09257_),
    .X(_09258_));
 sky130_fd_sc_hd__inv_2 _16697_ (.A(_09258_),
    .Y(_09259_));
 sky130_fd_sc_hd__or3_1 _16698_ (.A(_09247_),
    .B(_09240_),
    .C(_09257_),
    .X(_09260_));
 sky130_fd_sc_hd__nand2_1 _16699_ (.A(_09259_),
    .B(_09260_),
    .Y(_09261_));
 sky130_fd_sc_hd__or2_2 _16700_ (.A(_09243_),
    .B(_09261_),
    .X(_09262_));
 sky130_fd_sc_hd__a21oi_1 _16701_ (.A1(_09243_),
    .A2(_09261_),
    .B1(_05399_),
    .Y(_09263_));
 sky130_fd_sc_hd__a22o_1 _16702_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[3] ),
    .A2(_08066_),
    .B1(_09262_),
    .B2(_09263_),
    .X(_09264_));
 sky130_fd_sc_hd__and2_1 _16703_ (.A(_08831_),
    .B(_09264_),
    .X(_09265_));
 sky130_fd_sc_hd__clkbuf_1 _16704_ (.A(_09265_),
    .X(_00560_));
 sky130_fd_sc_hd__buf_6 _16705_ (.A(_05787_),
    .X(_09266_));
 sky130_fd_sc_hd__nand2_1 _16706_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[2] ),
    .B(_09197_),
    .Y(_09267_));
 sky130_fd_sc_hd__nand4_4 _16707_ (.A(_09207_),
    .B(_09203_),
    .C(_09186_),
    .D(net1120),
    .Y(_09268_));
 sky130_fd_sc_hd__a22o_1 _16708_ (.A1(_09207_),
    .A2(_09186_),
    .B1(net1120),
    .B2(_09203_),
    .X(_09269_));
 sky130_fd_sc_hd__nand3b_2 _16709_ (.A_N(_09267_),
    .B(_09268_),
    .C(_09269_),
    .Y(_09270_));
 sky130_fd_sc_hd__a21bo_1 _16710_ (.A1(_09268_),
    .A2(_09269_),
    .B1_N(_09267_),
    .X(_09271_));
 sky130_fd_sc_hd__and2_1 _16711_ (.A(_09270_),
    .B(_09271_),
    .X(_09272_));
 sky130_fd_sc_hd__a21bo_1 _16712_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[3] ),
    .A2(_09248_),
    .B1_N(_09249_),
    .X(_09273_));
 sky130_fd_sc_hd__a22o_1 _16713_ (.A1(_09193_),
    .A2(_09202_),
    .B1(_09206_),
    .B2(_09188_),
    .X(_09274_));
 sky130_fd_sc_hd__nand4_1 _16714_ (.A(_09193_),
    .B(_09188_),
    .C(_09202_),
    .D(_09206_),
    .Y(_09275_));
 sky130_fd_sc_hd__and3_1 _16715_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[4] ),
    .B(_09274_),
    .C(_09275_),
    .X(_09276_));
 sky130_fd_sc_hd__a21oi_1 _16716_ (.A1(_09274_),
    .A2(_09275_),
    .B1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[4] ),
    .Y(_09277_));
 sky130_fd_sc_hd__or3_4 _16717_ (.A(_09255_),
    .B(_09276_),
    .C(_09277_),
    .X(_09278_));
 sky130_fd_sc_hd__o21ai_1 _16718_ (.A1(_09276_),
    .A2(_09277_),
    .B1(_09255_),
    .Y(_09279_));
 sky130_fd_sc_hd__nand3_2 _16719_ (.A(_09273_),
    .B(_09278_),
    .C(_09279_),
    .Y(_09280_));
 sky130_fd_sc_hd__a21o_1 _16720_ (.A1(_09278_),
    .A2(_09279_),
    .B1(_09273_),
    .X(_09281_));
 sky130_fd_sc_hd__nand3_4 _16721_ (.A(_09272_),
    .B(_09280_),
    .C(_09281_),
    .Y(_09282_));
 sky130_fd_sc_hd__a21o_1 _16722_ (.A1(_09280_),
    .A2(_09281_),
    .B1(_09272_),
    .X(_09283_));
 sky130_fd_sc_hd__inv_2 _16723_ (.A(_09256_),
    .Y(_09284_));
 sky130_fd_sc_hd__nand2_1 _16724_ (.A(_09251_),
    .B(_09252_),
    .Y(_09285_));
 sky130_fd_sc_hd__o21ai_1 _16725_ (.A1(_09253_),
    .A2(_09284_),
    .B1(_09285_),
    .Y(_09286_));
 sky130_fd_sc_hd__nand3_2 _16726_ (.A(_09282_),
    .B(_09283_),
    .C(_09286_),
    .Y(_09287_));
 sky130_fd_sc_hd__a21o_1 _16727_ (.A1(_09282_),
    .A2(_09283_),
    .B1(_09286_),
    .X(_09288_));
 sky130_fd_sc_hd__nand2_2 _16728_ (.A(_09287_),
    .B(_09288_),
    .Y(_09289_));
 sky130_fd_sc_hd__nand2_1 _16729_ (.A(_09259_),
    .B(_09262_),
    .Y(_09290_));
 sky130_fd_sc_hd__nor2_1 _16730_ (.A(_09289_),
    .B(_09290_),
    .Y(_09291_));
 sky130_fd_sc_hd__buf_8 _16731_ (.A(_05327_),
    .X(_09292_));
 sky130_fd_sc_hd__a21o_1 _16732_ (.A1(_09289_),
    .A2(_09290_),
    .B1(_09292_),
    .X(_09293_));
 sky130_fd_sc_hd__o221a_1 _16733_ (.A1(net1081),
    .A2(_09266_),
    .B1(_09291_),
    .B2(_09293_),
    .C1(_07708_),
    .X(_00561_));
 sky130_fd_sc_hd__nor2_1 _16734_ (.A(_09262_),
    .B(_09289_),
    .Y(_09294_));
 sky130_fd_sc_hd__a21bo_1 _16735_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[4] ),
    .A2(_09274_),
    .B1_N(_09275_),
    .X(_09295_));
 sky130_fd_sc_hd__a22o_1 _16736_ (.A1(_09193_),
    .A2(net216),
    .B1(_09209_),
    .B2(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[0] ),
    .X(_09296_));
 sky130_fd_sc_hd__nand4_2 _16737_ (.A(_09193_),
    .B(_09188_),
    .C(net217),
    .D(_09210_),
    .Y(_09297_));
 sky130_fd_sc_hd__and3_1 _16738_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[5] ),
    .B(_09296_),
    .C(_09297_),
    .X(_09298_));
 sky130_fd_sc_hd__a21oi_1 _16739_ (.A1(_09296_),
    .A2(_09297_),
    .B1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[5] ),
    .Y(_09299_));
 sky130_fd_sc_hd__a211o_1 _16740_ (.A1(_09268_),
    .A2(_09270_),
    .B1(_09298_),
    .C1(_09299_),
    .X(_09300_));
 sky130_fd_sc_hd__o211ai_2 _16741_ (.A1(_09298_),
    .A2(_09299_),
    .B1(_09268_),
    .C1(_09270_),
    .Y(_09301_));
 sky130_fd_sc_hd__nand3_2 _16742_ (.A(_09295_),
    .B(_09300_),
    .C(_09301_),
    .Y(_09302_));
 sky130_fd_sc_hd__a21o_1 _16743_ (.A1(_09300_),
    .A2(_09301_),
    .B1(_09295_),
    .X(_09303_));
 sky130_fd_sc_hd__a22o_1 _16744_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[4] ),
    .A2(net1119),
    .B1(net225),
    .B2(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[3] ),
    .X(_09304_));
 sky130_fd_sc_hd__nand4_4 _16745_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[3] ),
    .C(net1119),
    .D(net225),
    .Y(_09305_));
 sky130_fd_sc_hd__nand4_2 _16746_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[2] ),
    .B(_09202_),
    .C(_09304_),
    .D(_09305_),
    .Y(_09306_));
 sky130_fd_sc_hd__a22o_1 _16747_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[2] ),
    .A2(_09202_),
    .B1(_09304_),
    .B2(_09305_),
    .X(_09307_));
 sky130_fd_sc_hd__and4_1 _16748_ (.A(_09211_),
    .B(_09187_),
    .C(_09306_),
    .D(_09307_),
    .X(_09308_));
 sky130_fd_sc_hd__a22oi_1 _16749_ (.A1(_09211_),
    .A2(_09187_),
    .B1(_09306_),
    .B2(_09307_),
    .Y(_09309_));
 sky130_fd_sc_hd__nor2_1 _16750_ (.A(_09308_),
    .B(_09309_),
    .Y(_09310_));
 sky130_fd_sc_hd__and3_1 _16751_ (.A(_09302_),
    .B(_09303_),
    .C(_09310_),
    .X(_09311_));
 sky130_fd_sc_hd__a21oi_1 _16752_ (.A1(_09302_),
    .A2(_09303_),
    .B1(_09310_),
    .Y(_09312_));
 sky130_fd_sc_hd__nor3_2 _16753_ (.A(_09282_),
    .B(_09311_),
    .C(_09312_),
    .Y(_09313_));
 sky130_fd_sc_hd__o21a_1 _16754_ (.A1(_09311_),
    .A2(_09312_),
    .B1(_09282_),
    .X(_09314_));
 sky130_fd_sc_hd__nand2_1 _16755_ (.A(_09278_),
    .B(_09280_),
    .Y(_09315_));
 sky130_fd_sc_hd__nor3b_1 _16756_ (.A(net170),
    .B(_09314_),
    .C_N(_09315_),
    .Y(_09316_));
 sky130_fd_sc_hd__o21ba_1 _16757_ (.A1(_09313_),
    .A2(_09314_),
    .B1_N(_09315_),
    .X(_09317_));
 sky130_fd_sc_hd__or2_4 _16758_ (.A(_09316_),
    .B(_09317_),
    .X(_09318_));
 sky130_fd_sc_hd__o21a_1 _16759_ (.A1(_09259_),
    .A2(_09289_),
    .B1(_09287_),
    .X(_09319_));
 sky130_fd_sc_hd__xnor2_2 _16760_ (.A(_09318_),
    .B(_09319_),
    .Y(_09320_));
 sky130_fd_sc_hd__xnor2_1 _16761_ (.A(_09294_),
    .B(_09320_),
    .Y(_09321_));
 sky130_fd_sc_hd__mux2_1 _16762_ (.A0(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[5] ),
    .A1(_09321_),
    .S(_08307_),
    .X(_09322_));
 sky130_fd_sc_hd__and2_1 _16763_ (.A(_08831_),
    .B(_09322_),
    .X(_09323_));
 sky130_fd_sc_hd__clkbuf_1 _16764_ (.A(_09323_),
    .X(_00562_));
 sky130_fd_sc_hd__a21bo_1 _16765_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[5] ),
    .A2(_09296_),
    .B1_N(_09297_),
    .X(_09324_));
 sky130_fd_sc_hd__a22o_1 _16766_ (.A1(_09193_),
    .A2(_09209_),
    .B1(_09214_),
    .B2(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[0] ),
    .X(_09325_));
 sky130_fd_sc_hd__nand4_1 _16767_ (.A(_09193_),
    .B(_09188_),
    .C(_09210_),
    .D(net202),
    .Y(_09326_));
 sky130_fd_sc_hd__and3_1 _16768_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[6] ),
    .B(_09325_),
    .C(_09326_),
    .X(_09327_));
 sky130_fd_sc_hd__a21oi_1 _16769_ (.A1(_09325_),
    .A2(_09326_),
    .B1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[6] ),
    .Y(_09328_));
 sky130_fd_sc_hd__a211o_4 _16770_ (.A1(_09305_),
    .A2(_09306_),
    .B1(_09327_),
    .C1(_09328_),
    .X(_09329_));
 sky130_fd_sc_hd__o211ai_2 _16771_ (.A1(_09327_),
    .A2(_09328_),
    .B1(_09305_),
    .C1(_09306_),
    .Y(_09330_));
 sky130_fd_sc_hd__nand3_2 _16772_ (.A(_09324_),
    .B(_09329_),
    .C(_09330_),
    .Y(_09331_));
 sky130_fd_sc_hd__a21o_1 _16773_ (.A1(_09329_),
    .A2(_09330_),
    .B1(_09324_),
    .X(_09332_));
 sky130_fd_sc_hd__a22o_1 _16774_ (.A1(_09207_),
    .A2(_09197_),
    .B1(_09201_),
    .B2(_09203_),
    .X(_09333_));
 sky130_fd_sc_hd__nand4_2 _16775_ (.A(_09207_),
    .B(_09203_),
    .C(_09197_),
    .D(_09202_),
    .Y(_09334_));
 sky130_fd_sc_hd__nand4_2 _16776_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[2] ),
    .B(_09206_),
    .C(_09333_),
    .D(_09334_),
    .Y(_09335_));
 sky130_fd_sc_hd__a22o_1 _16777_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[2] ),
    .A2(_09206_),
    .B1(_09333_),
    .B2(_09334_),
    .X(_09336_));
 sky130_fd_sc_hd__a22oi_1 _16778_ (.A1(_09213_),
    .A2(_09186_),
    .B1(_09192_),
    .B2(_09211_),
    .Y(_09337_));
 sky130_fd_sc_hd__and4_1 _16779_ (.A(_09213_),
    .B(_09211_),
    .C(_09186_),
    .D(_09192_),
    .X(_09338_));
 sky130_fd_sc_hd__nor2_1 _16780_ (.A(_09337_),
    .B(_09338_),
    .Y(_09339_));
 sky130_fd_sc_hd__nand3_1 _16781_ (.A(_09335_),
    .B(_09336_),
    .C(_09339_),
    .Y(_09340_));
 sky130_fd_sc_hd__a21o_1 _16782_ (.A1(_09335_),
    .A2(_09336_),
    .B1(_09339_),
    .X(_09341_));
 sky130_fd_sc_hd__nand3_2 _16783_ (.A(_09308_),
    .B(_09340_),
    .C(_09341_),
    .Y(_09342_));
 sky130_fd_sc_hd__a21o_1 _16784_ (.A1(_09340_),
    .A2(_09341_),
    .B1(_09308_),
    .X(_09343_));
 sky130_fd_sc_hd__nand4_2 _16785_ (.A(_09331_),
    .B(_09332_),
    .C(_09342_),
    .D(_09343_),
    .Y(_09344_));
 sky130_fd_sc_hd__a22o_1 _16786_ (.A1(_09331_),
    .A2(_09332_),
    .B1(_09342_),
    .B2(_09343_),
    .X(_09345_));
 sky130_fd_sc_hd__and3_1 _16787_ (.A(_09311_),
    .B(_09344_),
    .C(_09345_),
    .X(_09346_));
 sky130_fd_sc_hd__a21oi_1 _16788_ (.A1(_09344_),
    .A2(_09345_),
    .B1(_09311_),
    .Y(_09347_));
 sky130_fd_sc_hd__a211o_1 _16789_ (.A1(_09300_),
    .A2(_09302_),
    .B1(_09346_),
    .C1(_09347_),
    .X(_09348_));
 sky130_fd_sc_hd__o211ai_1 _16790_ (.A1(_09346_),
    .A2(_09347_),
    .B1(_09300_),
    .C1(_09302_),
    .Y(_09349_));
 sky130_fd_sc_hd__o211a_1 _16791_ (.A1(net170),
    .A2(_09316_),
    .B1(_09348_),
    .C1(_09349_),
    .X(_09350_));
 sky130_fd_sc_hd__a211oi_1 _16792_ (.A1(_09348_),
    .A2(_09349_),
    .B1(net170),
    .C1(_09316_),
    .Y(_09351_));
 sky130_fd_sc_hd__or4_1 _16793_ (.A(_09287_),
    .B(_09318_),
    .C(_09350_),
    .D(_09351_),
    .X(_09352_));
 sky130_fd_sc_hd__o22ai_1 _16794_ (.A1(_09287_),
    .A2(_09318_),
    .B1(_09350_),
    .B2(_09351_),
    .Y(_09353_));
 sky130_fd_sc_hd__and2_1 _16795_ (.A(_09352_),
    .B(_09353_),
    .X(_09354_));
 sky130_fd_sc_hd__or2_1 _16796_ (.A(_09259_),
    .B(_09289_),
    .X(_09355_));
 sky130_fd_sc_hd__o32ai_4 _16797_ (.A1(_09262_),
    .A2(_09289_),
    .A3(_09320_),
    .B1(_09355_),
    .B2(_09318_),
    .Y(_09356_));
 sky130_fd_sc_hd__xor2_1 _16798_ (.A(_09354_),
    .B(_09356_),
    .X(_09357_));
 sky130_fd_sc_hd__mux2_1 _16799_ (.A0(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[6] ),
    .A1(_09357_),
    .S(_08307_),
    .X(_09358_));
 sky130_fd_sc_hd__and2_1 _16800_ (.A(_08831_),
    .B(_09358_),
    .X(_09359_));
 sky130_fd_sc_hd__clkbuf_1 _16801_ (.A(_09359_),
    .X(_00563_));
 sky130_fd_sc_hd__inv_2 _16802_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[7] ),
    .Y(_09360_));
 sky130_fd_sc_hd__buf_2 _16803_ (.A(_09360_),
    .X(_09361_));
 sky130_fd_sc_hd__a21boi_1 _16804_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[6] ),
    .A2(_09325_),
    .B1_N(_09326_),
    .Y(_09362_));
 sky130_fd_sc_hd__nand2_1 _16805_ (.A(_09334_),
    .B(_09335_),
    .Y(_09363_));
 sky130_fd_sc_hd__a22o_1 _16806_ (.A1(_09193_),
    .A2(_09215_),
    .B1(_09218_),
    .B2(_09188_),
    .X(_09364_));
 sky130_fd_sc_hd__nand4_1 _16807_ (.A(_09193_),
    .B(_09188_),
    .C(_09215_),
    .D(net219),
    .Y(_09365_));
 sky130_fd_sc_hd__nand2_1 _16808_ (.A(_09364_),
    .B(_09365_),
    .Y(_09366_));
 sky130_fd_sc_hd__xor2_1 _16809_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[7] ),
    .B(_09366_),
    .X(_09367_));
 sky130_fd_sc_hd__xnor2_1 _16810_ (.A(_09363_),
    .B(_09367_),
    .Y(_09368_));
 sky130_fd_sc_hd__xnor2_1 _16811_ (.A(_09362_),
    .B(_09368_),
    .Y(_09369_));
 sky130_fd_sc_hd__and3_1 _16812_ (.A(_09335_),
    .B(_09336_),
    .C(_09339_),
    .X(_09370_));
 sky130_fd_sc_hd__nand2_1 _16813_ (.A(_09198_),
    .B(_09210_),
    .Y(_09371_));
 sky130_fd_sc_hd__a22oi_1 _16814_ (.A1(_09207_),
    .A2(_09202_),
    .B1(_09206_),
    .B2(_09203_),
    .Y(_09372_));
 sky130_fd_sc_hd__and4_1 _16815_ (.A(_09207_),
    .B(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[3] ),
    .C(_09201_),
    .D(_09206_),
    .X(_09373_));
 sky130_fd_sc_hd__nor2_1 _16816_ (.A(_09372_),
    .B(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__xnor2_1 _16817_ (.A(_09371_),
    .B(_09374_),
    .Y(_09375_));
 sky130_fd_sc_hd__and2_1 _16818_ (.A(_09211_),
    .B(_09197_),
    .X(_09376_));
 sky130_fd_sc_hd__inv_2 _16819_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[6] ),
    .Y(_09377_));
 sky130_fd_sc_hd__or4b_4 _16820_ (.A(_09360_),
    .B(_09377_),
    .C(_09186_),
    .D_N(_09191_),
    .X(_09378_));
 sky130_fd_sc_hd__a2bb2o_1 _16821_ (.A1_N(_09361_),
    .A2_N(_09186_),
    .B1(_09191_),
    .B2(_09213_),
    .X(_09379_));
 sky130_fd_sc_hd__nand3_1 _16822_ (.A(_09376_),
    .B(_09378_),
    .C(_09379_),
    .Y(_09380_));
 sky130_fd_sc_hd__a21o_1 _16823_ (.A1(_09378_),
    .A2(_09379_),
    .B1(_09376_),
    .X(_09381_));
 sky130_fd_sc_hd__nand3_1 _16824_ (.A(_09338_),
    .B(_09380_),
    .C(_09381_),
    .Y(_09382_));
 sky130_fd_sc_hd__a21o_1 _16825_ (.A1(_09380_),
    .A2(_09381_),
    .B1(_09338_),
    .X(_09383_));
 sky130_fd_sc_hd__nand3_1 _16826_ (.A(_09375_),
    .B(_09382_),
    .C(_09383_),
    .Y(_09384_));
 sky130_fd_sc_hd__a21o_1 _16827_ (.A1(_09382_),
    .A2(_09383_),
    .B1(_09375_),
    .X(_09385_));
 sky130_fd_sc_hd__nand3_2 _16828_ (.A(_09370_),
    .B(_09384_),
    .C(_09385_),
    .Y(_09386_));
 sky130_fd_sc_hd__a21o_1 _16829_ (.A1(_09384_),
    .A2(_09385_),
    .B1(_09370_),
    .X(_09387_));
 sky130_fd_sc_hd__nand3_2 _16830_ (.A(_09369_),
    .B(_09386_),
    .C(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__a21o_1 _16831_ (.A1(_09386_),
    .A2(_09387_),
    .B1(_09369_),
    .X(_09389_));
 sky130_fd_sc_hd__nand2_1 _16832_ (.A(_09342_),
    .B(_09344_),
    .Y(_09390_));
 sky130_fd_sc_hd__and3_1 _16833_ (.A(_09388_),
    .B(_09389_),
    .C(_09390_),
    .X(_09391_));
 sky130_fd_sc_hd__a21oi_1 _16834_ (.A1(_09388_),
    .A2(_09389_),
    .B1(_09390_),
    .Y(_09392_));
 sky130_fd_sc_hd__a211oi_4 _16835_ (.A1(_09329_),
    .A2(_09331_),
    .B1(_09391_),
    .C1(_09392_),
    .Y(_09393_));
 sky130_fd_sc_hd__o211a_1 _16836_ (.A1(_09391_),
    .A2(_09392_),
    .B1(_09329_),
    .C1(_09331_),
    .X(_09394_));
 sky130_fd_sc_hd__and2b_1 _16837_ (.A_N(_09346_),
    .B(_09348_),
    .X(_09395_));
 sky130_fd_sc_hd__nor3_2 _16838_ (.A(_09393_),
    .B(_09394_),
    .C(_09395_),
    .Y(_09396_));
 sky130_fd_sc_hd__o21ai_1 _16839_ (.A1(_09393_),
    .A2(_09394_),
    .B1(_09395_),
    .Y(_09397_));
 sky130_fd_sc_hd__or3b_1 _16840_ (.A(_09361_),
    .B(_09396_),
    .C_N(_09397_),
    .X(_09398_));
 sky130_fd_sc_hd__or3_1 _16841_ (.A(_09393_),
    .B(_09394_),
    .C(_09395_),
    .X(_09399_));
 sky130_fd_sc_hd__a21o_1 _16842_ (.A1(_09399_),
    .A2(_09397_),
    .B1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[7] ),
    .X(_09400_));
 sky130_fd_sc_hd__and3_1 _16843_ (.A(_09350_),
    .B(_09398_),
    .C(_09400_),
    .X(_09401_));
 sky130_fd_sc_hd__a21o_1 _16844_ (.A1(_09398_),
    .A2(_09400_),
    .B1(_09350_),
    .X(_09402_));
 sky130_fd_sc_hd__and2b_1 _16845_ (.A_N(_09401_),
    .B(_09402_),
    .X(_09403_));
 sky130_fd_sc_hd__a21bo_1 _16846_ (.A1(_09354_),
    .A2(_09356_),
    .B1_N(_09352_),
    .X(_09404_));
 sky130_fd_sc_hd__or2_1 _16847_ (.A(_09403_),
    .B(_09404_),
    .X(_09405_));
 sky130_fd_sc_hd__a21oi_1 _16848_ (.A1(_09403_),
    .A2(_09404_),
    .B1(_05399_),
    .Y(_09406_));
 sky130_fd_sc_hd__a22o_1 _16849_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[7] ),
    .A2(_08066_),
    .B1(_09405_),
    .B2(_09406_),
    .X(_09407_));
 sky130_fd_sc_hd__and2_1 _16850_ (.A(_08831_),
    .B(_09407_),
    .X(_09408_));
 sky130_fd_sc_hd__clkbuf_1 _16851_ (.A(_09408_),
    .X(_00564_));
 sky130_fd_sc_hd__a21oi_4 _16852_ (.A1(_09402_),
    .A2(_09404_),
    .B1(_09401_),
    .Y(_09409_));
 sky130_fd_sc_hd__nor2_2 _16853_ (.A(_09391_),
    .B(_09393_),
    .Y(_09410_));
 sky130_fd_sc_hd__or2b_1 _16854_ (.A(_09367_),
    .B_N(_09363_),
    .X(_09411_));
 sky130_fd_sc_hd__or2b_1 _16855_ (.A(_09362_),
    .B_N(_09368_),
    .X(_09412_));
 sky130_fd_sc_hd__nand2_1 _16856_ (.A(_09411_),
    .B(_09412_),
    .Y(_09413_));
 sky130_fd_sc_hd__a21boi_1 _16857_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[7] ),
    .A2(_09364_),
    .B1_N(_09365_),
    .Y(_09414_));
 sky130_fd_sc_hd__a31o_1 _16858_ (.A1(_09198_),
    .A2(_09210_),
    .A3(_09374_),
    .B1(_09373_),
    .X(_09415_));
 sky130_fd_sc_hd__and3_1 _16859_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[1] ),
    .B(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[0] ),
    .C(_09217_),
    .X(_09416_));
 sky130_fd_sc_hd__clkbuf_4 _16860_ (.A(_09416_),
    .X(_09417_));
 sky130_fd_sc_hd__o21ai_4 _16861_ (.A1(_09193_),
    .A2(_09188_),
    .B1(net219),
    .Y(_09418_));
 sky130_fd_sc_hd__nor2_8 _16862_ (.A(_09418_),
    .B(_09417_),
    .Y(_09419_));
 sky130_fd_sc_hd__xnor2_1 _16863_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[8] ),
    .B(_09419_),
    .Y(_09420_));
 sky130_fd_sc_hd__xnor2_1 _16864_ (.A(_09415_),
    .B(_09420_),
    .Y(_09421_));
 sky130_fd_sc_hd__xnor2_1 _16865_ (.A(_09414_),
    .B(_09421_),
    .Y(_09422_));
 sky130_fd_sc_hd__nand2_1 _16866_ (.A(_09198_),
    .B(_09215_),
    .Y(_09423_));
 sky130_fd_sc_hd__a22oi_1 _16867_ (.A1(_09207_),
    .A2(_09206_),
    .B1(_09210_),
    .B2(_09203_),
    .Y(_09424_));
 sky130_fd_sc_hd__and4_1 _16868_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[3] ),
    .C(net215),
    .D(_09209_),
    .X(_09425_));
 sky130_fd_sc_hd__nor2_1 _16869_ (.A(_09424_),
    .B(_09425_),
    .Y(_09426_));
 sky130_fd_sc_hd__xnor2_1 _16870_ (.A(_09423_),
    .B(_09426_),
    .Y(_09427_));
 sky130_fd_sc_hd__and2_1 _16871_ (.A(_09211_),
    .B(_09201_),
    .X(_09428_));
 sky130_fd_sc_hd__or4b_4 _16872_ (.A(_09360_),
    .B(_09377_),
    .C(_09191_),
    .D_N(_09196_),
    .X(_09429_));
 sky130_fd_sc_hd__a2bb2o_1 _16873_ (.A1_N(_09361_),
    .A2_N(_09191_),
    .B1(net224),
    .B2(_09213_),
    .X(_09430_));
 sky130_fd_sc_hd__nand3_1 _16874_ (.A(_09428_),
    .B(_09429_),
    .C(_09430_),
    .Y(_09431_));
 sky130_fd_sc_hd__a21o_1 _16875_ (.A1(_09429_),
    .A2(_09430_),
    .B1(_09428_),
    .X(_09432_));
 sky130_fd_sc_hd__a21bo_1 _16876_ (.A1(_09376_),
    .A2(_09379_),
    .B1_N(_09378_),
    .X(_09433_));
 sky130_fd_sc_hd__nand3_1 _16877_ (.A(_09431_),
    .B(_09432_),
    .C(_09433_),
    .Y(_09434_));
 sky130_fd_sc_hd__a21o_1 _16878_ (.A1(_09431_),
    .A2(_09432_),
    .B1(_09433_),
    .X(_09435_));
 sky130_fd_sc_hd__nand3_1 _16879_ (.A(_09427_),
    .B(_09434_),
    .C(_09435_),
    .Y(_09436_));
 sky130_fd_sc_hd__a21o_1 _16880_ (.A1(_09434_),
    .A2(_09435_),
    .B1(_09427_),
    .X(_09437_));
 sky130_fd_sc_hd__a21bo_1 _16881_ (.A1(_09375_),
    .A2(_09383_),
    .B1_N(_09382_),
    .X(_09438_));
 sky130_fd_sc_hd__nand3_2 _16882_ (.A(_09436_),
    .B(_09437_),
    .C(_09438_),
    .Y(_09439_));
 sky130_fd_sc_hd__a21o_1 _16883_ (.A1(_09436_),
    .A2(_09437_),
    .B1(_09438_),
    .X(_09440_));
 sky130_fd_sc_hd__and3_1 _16884_ (.A(_09422_),
    .B(_09439_),
    .C(_09440_),
    .X(_09441_));
 sky130_fd_sc_hd__a21oi_1 _16885_ (.A1(_09439_),
    .A2(_09440_),
    .B1(_09422_),
    .Y(_09442_));
 sky130_fd_sc_hd__a211oi_2 _16886_ (.A1(_09386_),
    .A2(_09388_),
    .B1(_09441_),
    .C1(_09442_),
    .Y(_09443_));
 sky130_fd_sc_hd__o211a_1 _16887_ (.A1(_09441_),
    .A2(_09442_),
    .B1(_09386_),
    .C1(_09388_),
    .X(_09444_));
 sky130_fd_sc_hd__nor2_1 _16888_ (.A(_09443_),
    .B(_09444_),
    .Y(_09445_));
 sky130_fd_sc_hd__xor2_1 _16889_ (.A(_09413_),
    .B(_09445_),
    .X(_09446_));
 sky130_fd_sc_hd__xnor2_2 _16890_ (.A(_09410_),
    .B(net183),
    .Y(_09447_));
 sky130_fd_sc_hd__a21o_1 _16891_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[7] ),
    .A2(_09397_),
    .B1(_09396_),
    .X(_09448_));
 sky130_fd_sc_hd__xnor2_2 _16892_ (.A(_09447_),
    .B(_09448_),
    .Y(_09449_));
 sky130_fd_sc_hd__xor2_1 _16893_ (.A(_09409_),
    .B(_09449_),
    .X(_09450_));
 sky130_fd_sc_hd__or2_1 _16894_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[8] ),
    .B(_07866_),
    .X(_09451_));
 sky130_fd_sc_hd__o211a_1 _16895_ (.A1(_08870_),
    .A2(_09450_),
    .B1(_09451_),
    .C1(_09231_),
    .X(_00565_));
 sky130_fd_sc_hd__nand2_1 _16896_ (.A(_09447_),
    .B(_09448_),
    .Y(_09452_));
 sky130_fd_sc_hd__o21ai_1 _16897_ (.A1(_09409_),
    .A2(_09449_),
    .B1(_09452_),
    .Y(_09453_));
 sky130_fd_sc_hd__or2b_1 _16898_ (.A(_09410_),
    .B_N(_09446_),
    .X(_09454_));
 sky130_fd_sc_hd__or2b_1 _16899_ (.A(_09420_),
    .B_N(_09415_),
    .X(_09455_));
 sky130_fd_sc_hd__or2b_1 _16900_ (.A(_09414_),
    .B_N(_09421_),
    .X(_09456_));
 sky130_fd_sc_hd__nand2_1 _16901_ (.A(_09455_),
    .B(_09456_),
    .Y(_09457_));
 sky130_fd_sc_hd__nand3_1 _16902_ (.A(_09422_),
    .B(_09439_),
    .C(_09440_),
    .Y(_09458_));
 sky130_fd_sc_hd__o21a_2 _16903_ (.A1(_09194_),
    .A2(_09189_),
    .B1(_09219_),
    .X(_09459_));
 sky130_fd_sc_hd__a21o_1 _16904_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[8] ),
    .A2(_09459_),
    .B1(_09417_),
    .X(_09460_));
 sky130_fd_sc_hd__a31o_1 _16905_ (.A1(_09198_),
    .A2(_09215_),
    .A3(_09426_),
    .B1(_09425_),
    .X(_09461_));
 sky130_fd_sc_hd__xnor2_1 _16906_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[9] ),
    .B(_09419_),
    .Y(_09462_));
 sky130_fd_sc_hd__xnor2_1 _16907_ (.A(_09461_),
    .B(_09462_),
    .Y(_09463_));
 sky130_fd_sc_hd__xor2_1 _16908_ (.A(_09460_),
    .B(_09463_),
    .X(_09464_));
 sky130_fd_sc_hd__nand2_2 _16909_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[2] ),
    .B(_09218_),
    .Y(_09465_));
 sky130_fd_sc_hd__and3_1 _16910_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[3] ),
    .C(_09210_),
    .X(_09466_));
 sky130_fd_sc_hd__a22o_1 _16911_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[4] ),
    .A2(_09209_),
    .B1(net203),
    .B2(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[3] ),
    .X(_09467_));
 sky130_fd_sc_hd__a21bo_1 _16912_ (.A1(_09215_),
    .A2(_09466_),
    .B1_N(_09467_),
    .X(_09468_));
 sky130_fd_sc_hd__xor2_1 _16913_ (.A(_09465_),
    .B(_09468_),
    .X(_09469_));
 sky130_fd_sc_hd__and2_1 _16914_ (.A(_09211_),
    .B(_09206_),
    .X(_09470_));
 sky130_fd_sc_hd__or4b_4 _16915_ (.A(_09360_),
    .B(_09377_),
    .C(_09196_),
    .D_N(_09201_),
    .X(_09471_));
 sky130_fd_sc_hd__a2bb2o_1 _16916_ (.A1_N(_09361_),
    .A2_N(net223),
    .B1(_09201_),
    .B2(_09213_),
    .X(_09472_));
 sky130_fd_sc_hd__nand3_1 _16917_ (.A(_09470_),
    .B(_09471_),
    .C(_09472_),
    .Y(_09473_));
 sky130_fd_sc_hd__a21o_1 _16918_ (.A1(_09471_),
    .A2(_09472_),
    .B1(_09470_),
    .X(_09474_));
 sky130_fd_sc_hd__a21bo_1 _16919_ (.A1(_09428_),
    .A2(_09430_),
    .B1_N(_09429_),
    .X(_09475_));
 sky130_fd_sc_hd__nand3_1 _16920_ (.A(_09473_),
    .B(_09474_),
    .C(_09475_),
    .Y(_09476_));
 sky130_fd_sc_hd__a21o_1 _16921_ (.A1(_09473_),
    .A2(_09474_),
    .B1(_09475_),
    .X(_09477_));
 sky130_fd_sc_hd__nand3_1 _16922_ (.A(_09469_),
    .B(_09476_),
    .C(_09477_),
    .Y(_09478_));
 sky130_fd_sc_hd__a21o_1 _16923_ (.A1(_09476_),
    .A2(_09477_),
    .B1(_09469_),
    .X(_09479_));
 sky130_fd_sc_hd__a21bo_1 _16924_ (.A1(_09427_),
    .A2(_09435_),
    .B1_N(_09434_),
    .X(_09480_));
 sky130_fd_sc_hd__nand3_2 _16925_ (.A(_09478_),
    .B(_09479_),
    .C(_09480_),
    .Y(_09481_));
 sky130_fd_sc_hd__a21o_1 _16926_ (.A1(_09478_),
    .A2(_09479_),
    .B1(_09480_),
    .X(_09482_));
 sky130_fd_sc_hd__and3_1 _16927_ (.A(net200),
    .B(_09481_),
    .C(_09482_),
    .X(_09483_));
 sky130_fd_sc_hd__a21oi_1 _16928_ (.A1(_09481_),
    .A2(_09482_),
    .B1(net200),
    .Y(_09484_));
 sky130_fd_sc_hd__a211o_1 _16929_ (.A1(_09439_),
    .A2(_09458_),
    .B1(_09483_),
    .C1(_09484_),
    .X(_09485_));
 sky130_fd_sc_hd__o211ai_1 _16930_ (.A1(_09483_),
    .A2(_09484_),
    .B1(_09439_),
    .C1(_09458_),
    .Y(_09486_));
 sky130_fd_sc_hd__nand3_1 _16931_ (.A(_09457_),
    .B(_09485_),
    .C(_09486_),
    .Y(_09487_));
 sky130_fd_sc_hd__a21o_1 _16932_ (.A1(_09485_),
    .A2(_09486_),
    .B1(_09457_),
    .X(_09488_));
 sky130_fd_sc_hd__and2_1 _16933_ (.A(_09487_),
    .B(_09488_),
    .X(_09489_));
 sky130_fd_sc_hd__a21o_1 _16934_ (.A1(_09413_),
    .A2(_09445_),
    .B1(_09443_),
    .X(_09490_));
 sky130_fd_sc_hd__xnor2_2 _16935_ (.A(_09489_),
    .B(_09490_),
    .Y(_09491_));
 sky130_fd_sc_hd__xnor2_2 _16936_ (.A(_09454_),
    .B(_09491_),
    .Y(_09492_));
 sky130_fd_sc_hd__xnor2_1 _16937_ (.A(_09453_),
    .B(_09492_),
    .Y(_09493_));
 sky130_fd_sc_hd__clkbuf_8 _16938_ (.A(_05312_),
    .X(_09494_));
 sky130_fd_sc_hd__or2_1 _16939_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[9] ),
    .B(_09494_),
    .X(_09495_));
 sky130_fd_sc_hd__o211a_1 _16940_ (.A1(_08870_),
    .A2(_09493_),
    .B1(_09495_),
    .C1(_09231_),
    .X(_00566_));
 sky130_fd_sc_hd__buf_8 _16941_ (.A(_05326_),
    .X(_09496_));
 sky130_fd_sc_hd__nand2_1 _16942_ (.A(_09489_),
    .B(_09490_),
    .Y(_09497_));
 sky130_fd_sc_hd__and2b_1 _16943_ (.A_N(_09462_),
    .B(_09461_),
    .X(_09498_));
 sky130_fd_sc_hd__a21o_1 _16944_ (.A1(_09460_),
    .A2(_09463_),
    .B1(_09498_),
    .X(_09499_));
 sky130_fd_sc_hd__nand3_2 _16945_ (.A(_09464_),
    .B(_09481_),
    .C(_09482_),
    .Y(_09500_));
 sky130_fd_sc_hd__a21o_1 _16946_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[9] ),
    .A2(_09459_),
    .B1(_09417_),
    .X(_09501_));
 sky130_fd_sc_hd__a32o_1 _16947_ (.A1(_09198_),
    .A2(_09219_),
    .A3(_09467_),
    .B1(_09466_),
    .B2(_09215_),
    .X(_09502_));
 sky130_fd_sc_hd__xnor2_1 _16948_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[10] ),
    .B(_09419_),
    .Y(_09503_));
 sky130_fd_sc_hd__xnor2_1 _16949_ (.A(_09502_),
    .B(_09503_),
    .Y(_09504_));
 sky130_fd_sc_hd__xor2_1 _16950_ (.A(_09501_),
    .B(_09504_),
    .X(_09505_));
 sky130_fd_sc_hd__and3_1 _16951_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[3] ),
    .B(net203),
    .C(_09218_),
    .X(_09506_));
 sky130_fd_sc_hd__a22o_1 _16952_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[4] ),
    .A2(net203),
    .B1(_09218_),
    .B2(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[3] ),
    .X(_09507_));
 sky130_fd_sc_hd__a21bo_1 _16953_ (.A1(_09207_),
    .A2(_09506_),
    .B1_N(_09507_),
    .X(_09508_));
 sky130_fd_sc_hd__xor2_2 _16954_ (.A(_09465_),
    .B(_09508_),
    .X(_09509_));
 sky130_fd_sc_hd__and2_1 _16955_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[5] ),
    .B(_09209_),
    .X(_09510_));
 sky130_fd_sc_hd__or4b_4 _16956_ (.A(_09360_),
    .B(_09377_),
    .C(_09201_),
    .D_N(net227),
    .X(_09511_));
 sky130_fd_sc_hd__a2bb2o_2 _16957_ (.A1_N(_09360_),
    .A2_N(_09201_),
    .B1(net216),
    .B2(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[6] ),
    .X(_09512_));
 sky130_fd_sc_hd__nand3_1 _16958_ (.A(_09510_),
    .B(_09511_),
    .C(_09512_),
    .Y(_09513_));
 sky130_fd_sc_hd__a21o_1 _16959_ (.A1(_09511_),
    .A2(_09512_),
    .B1(_09510_),
    .X(_09514_));
 sky130_fd_sc_hd__a21bo_1 _16960_ (.A1(_09470_),
    .A2(_09472_),
    .B1_N(_09471_),
    .X(_09515_));
 sky130_fd_sc_hd__nand3_1 _16961_ (.A(_09513_),
    .B(net220),
    .C(_09515_),
    .Y(_09516_));
 sky130_fd_sc_hd__a21o_1 _16962_ (.A1(_09513_),
    .A2(_09514_),
    .B1(_09515_),
    .X(_09517_));
 sky130_fd_sc_hd__nand3_1 _16963_ (.A(_09509_),
    .B(_09516_),
    .C(net226),
    .Y(_09518_));
 sky130_fd_sc_hd__a21o_1 _16964_ (.A1(_09516_),
    .A2(_09517_),
    .B1(_09509_),
    .X(_09519_));
 sky130_fd_sc_hd__a21bo_2 _16965_ (.A1(_09469_),
    .A2(_09477_),
    .B1_N(_09476_),
    .X(_09520_));
 sky130_fd_sc_hd__nand3_4 _16966_ (.A(net204),
    .B(net201),
    .C(_09520_),
    .Y(_09521_));
 sky130_fd_sc_hd__a21o_1 _16967_ (.A1(_09518_),
    .A2(_09519_),
    .B1(_09520_),
    .X(_09522_));
 sky130_fd_sc_hd__and3_1 _16968_ (.A(_09505_),
    .B(_09521_),
    .C(_09522_),
    .X(_09523_));
 sky130_fd_sc_hd__a21oi_1 _16969_ (.A1(_09521_),
    .A2(_09522_),
    .B1(_09505_),
    .Y(_09524_));
 sky130_fd_sc_hd__a211o_1 _16970_ (.A1(_09481_),
    .A2(_09500_),
    .B1(_09523_),
    .C1(_09524_),
    .X(_09525_));
 sky130_fd_sc_hd__o211ai_2 _16971_ (.A1(_09523_),
    .A2(_09524_),
    .B1(_09481_),
    .C1(_09500_),
    .Y(_09526_));
 sky130_fd_sc_hd__and3_1 _16972_ (.A(_09499_),
    .B(_09525_),
    .C(_09526_),
    .X(_09527_));
 sky130_fd_sc_hd__a21oi_1 _16973_ (.A1(_09525_),
    .A2(_09526_),
    .B1(_09499_),
    .Y(_09528_));
 sky130_fd_sc_hd__a211oi_2 _16974_ (.A1(_09485_),
    .A2(_09487_),
    .B1(_09527_),
    .C1(_09528_),
    .Y(_09529_));
 sky130_fd_sc_hd__o211a_1 _16975_ (.A1(_09527_),
    .A2(_09528_),
    .B1(_09485_),
    .C1(_09487_),
    .X(_09530_));
 sky130_fd_sc_hd__or2_4 _16976_ (.A(_09529_),
    .B(_09530_),
    .X(_09531_));
 sky130_fd_sc_hd__xnor2_2 _16977_ (.A(_09497_),
    .B(_09531_),
    .Y(_09532_));
 sky130_fd_sc_hd__a21o_1 _16978_ (.A1(_09454_),
    .A2(_09452_),
    .B1(_09491_),
    .X(_09533_));
 sky130_fd_sc_hd__o31ai_1 _16979_ (.A1(_09409_),
    .A2(_09449_),
    .A3(_09492_),
    .B1(_09533_),
    .Y(_09534_));
 sky130_fd_sc_hd__or2b_1 _16980_ (.A(_09532_),
    .B_N(_09534_),
    .X(_09535_));
 sky130_fd_sc_hd__and2b_1 _16981_ (.A_N(_09534_),
    .B(_09532_),
    .X(_09536_));
 sky130_fd_sc_hd__nor2_1 _16982_ (.A(_05399_),
    .B(_09536_),
    .Y(_09537_));
 sky130_fd_sc_hd__a22o_1 _16983_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[10] ),
    .A2(_09496_),
    .B1(_09535_),
    .B2(_09537_),
    .X(_09538_));
 sky130_fd_sc_hd__and2_1 _16984_ (.A(_08831_),
    .B(_09538_),
    .X(_09539_));
 sky130_fd_sc_hd__clkbuf_1 _16985_ (.A(_09539_),
    .X(_00567_));
 sky130_fd_sc_hd__or2_1 _16986_ (.A(_09497_),
    .B(_09531_),
    .X(_09540_));
 sky130_fd_sc_hd__and2b_1 _16987_ (.A_N(_09503_),
    .B(_09502_),
    .X(_09541_));
 sky130_fd_sc_hd__a21o_1 _16988_ (.A1(_09501_),
    .A2(_09504_),
    .B1(_09541_),
    .X(_09542_));
 sky130_fd_sc_hd__nand3_1 _16989_ (.A(_09505_),
    .B(_09521_),
    .C(net214),
    .Y(_09543_));
 sky130_fd_sc_hd__a21o_1 _16990_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[10] ),
    .A2(_09459_),
    .B1(_09417_),
    .X(_09544_));
 sky130_fd_sc_hd__a32o_1 _16991_ (.A1(_09198_),
    .A2(_09219_),
    .A3(_09507_),
    .B1(_09506_),
    .B2(_09207_),
    .X(_09545_));
 sky130_fd_sc_hd__xnor2_1 _16992_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[11] ),
    .B(_09419_),
    .Y(_09546_));
 sky130_fd_sc_hd__xnor2_1 _16993_ (.A(_09545_),
    .B(_09546_),
    .Y(_09547_));
 sky130_fd_sc_hd__xor2_1 _16994_ (.A(_09544_),
    .B(_09547_),
    .X(_09548_));
 sky130_fd_sc_hd__and3_1 _16995_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[3] ),
    .C(_09217_),
    .X(_09549_));
 sky130_fd_sc_hd__o21ai_2 _16996_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[4] ),
    .A2(_09203_),
    .B1(_09218_),
    .Y(_09550_));
 sky130_fd_sc_hd__or3_4 _16997_ (.A(_09465_),
    .B(_09549_),
    .C(_09550_),
    .X(_09551_));
 sky130_fd_sc_hd__o21ai_4 _16998_ (.A1(_09549_),
    .A2(_09550_),
    .B1(_09465_),
    .Y(_09552_));
 sky130_fd_sc_hd__nand2_2 _16999_ (.A(_09551_),
    .B(_09552_),
    .Y(_09553_));
 sky130_fd_sc_hd__and2_1 _17000_ (.A(_09211_),
    .B(_09214_),
    .X(_09554_));
 sky130_fd_sc_hd__or4b_4 _17001_ (.A(_09360_),
    .B(_09377_),
    .C(_09205_),
    .D_N(_09209_),
    .X(_09555_));
 sky130_fd_sc_hd__a2bb2o_1 _17002_ (.A1_N(_09361_),
    .A2_N(_09205_),
    .B1(_09209_),
    .B2(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[6] ),
    .X(_09556_));
 sky130_fd_sc_hd__nand3_1 _17003_ (.A(_09554_),
    .B(net221),
    .C(_09556_),
    .Y(_09557_));
 sky130_fd_sc_hd__a21o_1 _17004_ (.A1(_09555_),
    .A2(_09556_),
    .B1(_09554_),
    .X(_09558_));
 sky130_fd_sc_hd__a21bo_1 _17005_ (.A1(_09510_),
    .A2(_09512_),
    .B1_N(_09511_),
    .X(_09559_));
 sky130_fd_sc_hd__and3_1 _17006_ (.A(_09557_),
    .B(_09558_),
    .C(_09559_),
    .X(_09560_));
 sky130_fd_sc_hd__a21oi_2 _17007_ (.A1(_09557_),
    .A2(_09558_),
    .B1(net1121),
    .Y(_09561_));
 sky130_fd_sc_hd__or3_4 _17008_ (.A(_09553_),
    .B(_09560_),
    .C(_09561_),
    .X(_09562_));
 sky130_fd_sc_hd__o21ai_2 _17009_ (.A1(net1117),
    .A2(_09561_),
    .B1(_09553_),
    .Y(_09563_));
 sky130_fd_sc_hd__a21bo_1 _17010_ (.A1(_09509_),
    .A2(net226),
    .B1_N(_09516_),
    .X(_09564_));
 sky130_fd_sc_hd__nand3_2 _17011_ (.A(_09562_),
    .B(_09563_),
    .C(_09564_),
    .Y(_09565_));
 sky130_fd_sc_hd__a21o_1 _17012_ (.A1(_09562_),
    .A2(_09563_),
    .B1(_09564_),
    .X(_09566_));
 sky130_fd_sc_hd__and3_1 _17013_ (.A(_09548_),
    .B(_09565_),
    .C(_09566_),
    .X(_09567_));
 sky130_fd_sc_hd__a21oi_1 _17014_ (.A1(_09565_),
    .A2(_09566_),
    .B1(_09548_),
    .Y(_09568_));
 sky130_fd_sc_hd__a211o_1 _17015_ (.A1(_09521_),
    .A2(_09543_),
    .B1(_09567_),
    .C1(_09568_),
    .X(_09569_));
 sky130_fd_sc_hd__o211ai_2 _17016_ (.A1(_09567_),
    .A2(_09568_),
    .B1(_09521_),
    .C1(_09543_),
    .Y(_09570_));
 sky130_fd_sc_hd__and3_1 _17017_ (.A(_09542_),
    .B(_09569_),
    .C(_09570_),
    .X(_09571_));
 sky130_fd_sc_hd__a21oi_1 _17018_ (.A1(_09569_),
    .A2(_09570_),
    .B1(_09542_),
    .Y(_09572_));
 sky130_fd_sc_hd__nor2_2 _17019_ (.A(_09571_),
    .B(_09572_),
    .Y(_09573_));
 sky130_fd_sc_hd__a21bo_1 _17020_ (.A1(_09499_),
    .A2(_09526_),
    .B1_N(_09525_),
    .X(_09574_));
 sky130_fd_sc_hd__xnor2_2 _17021_ (.A(_09573_),
    .B(_09574_),
    .Y(_09575_));
 sky130_fd_sc_hd__xnor2_2 _17022_ (.A(net1118),
    .B(_09575_),
    .Y(_09576_));
 sky130_fd_sc_hd__a21oi_1 _17023_ (.A1(_09540_),
    .A2(_09535_),
    .B1(_09576_),
    .Y(_09577_));
 sky130_fd_sc_hd__a31o_1 _17024_ (.A1(_09540_),
    .A2(_09535_),
    .A3(_09576_),
    .B1(_07439_),
    .X(_09578_));
 sky130_fd_sc_hd__o221a_1 _17025_ (.A1(net1040),
    .A2(_09266_),
    .B1(_09577_),
    .B2(_09578_),
    .C1(_07708_),
    .X(_00568_));
 sky130_fd_sc_hd__or2b_1 _17026_ (.A(_09532_),
    .B_N(_09576_),
    .X(_09579_));
 sky130_fd_sc_hd__or4b_4 _17027_ (.A(_09449_),
    .B(_09492_),
    .C(_09532_),
    .D_N(_09576_),
    .X(_09580_));
 sky130_fd_sc_hd__inv_2 _17028_ (.A(_09529_),
    .Y(_09581_));
 sky130_fd_sc_hd__a21o_1 _17029_ (.A1(_09581_),
    .A2(_09540_),
    .B1(_09575_),
    .X(_09582_));
 sky130_fd_sc_hd__o221a_4 _17030_ (.A1(_09533_),
    .A2(_09579_),
    .B1(_09580_),
    .B2(_09409_),
    .C1(_09582_),
    .X(_09583_));
 sky130_fd_sc_hd__nand2_1 _17031_ (.A(_09573_),
    .B(_09574_),
    .Y(_09584_));
 sky130_fd_sc_hd__a21bo_1 _17032_ (.A1(_09542_),
    .A2(_09570_),
    .B1_N(_09569_),
    .X(_09585_));
 sky130_fd_sc_hd__and2b_1 _17033_ (.A_N(_09546_),
    .B(_09545_),
    .X(_09586_));
 sky130_fd_sc_hd__a21o_1 _17034_ (.A1(_09544_),
    .A2(_09547_),
    .B1(_09586_),
    .X(_09587_));
 sky130_fd_sc_hd__nand3_2 _17035_ (.A(_09194_),
    .B(_09189_),
    .C(_09219_),
    .Y(_09588_));
 sky130_fd_sc_hd__nand2_1 _17036_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[11] ),
    .B(_09419_),
    .Y(_09589_));
 sky130_fd_sc_hd__nand2_1 _17037_ (.A(_09588_),
    .B(_09589_),
    .Y(_09590_));
 sky130_fd_sc_hd__o21ba_1 _17038_ (.A1(_09465_),
    .A2(_09550_),
    .B1_N(_09549_),
    .X(_09591_));
 sky130_fd_sc_hd__xnor2_1 _17039_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[12] ),
    .B(_09419_),
    .Y(_09592_));
 sky130_fd_sc_hd__xor2_1 _17040_ (.A(_09591_),
    .B(_09592_),
    .X(_09593_));
 sky130_fd_sc_hd__xor2_1 _17041_ (.A(_09590_),
    .B(_09593_),
    .X(_09594_));
 sky130_fd_sc_hd__a21bo_1 _17042_ (.A1(_09554_),
    .A2(_09556_),
    .B1_N(net222),
    .X(_09595_));
 sky130_fd_sc_hd__and2_1 _17043_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[5] ),
    .B(net219),
    .X(_09596_));
 sky130_fd_sc_hd__clkbuf_2 _17044_ (.A(_09596_),
    .X(_09597_));
 sky130_fd_sc_hd__or4b_4 _17045_ (.A(_09361_),
    .B(_09377_),
    .C(_09210_),
    .D_N(_09214_),
    .X(_09598_));
 sky130_fd_sc_hd__a2bb2o_1 _17046_ (.A1_N(_09361_),
    .A2_N(_09210_),
    .B1(net203),
    .B2(_09213_),
    .X(_09599_));
 sky130_fd_sc_hd__nand3_1 _17047_ (.A(_09597_),
    .B(_09598_),
    .C(_09599_),
    .Y(_09600_));
 sky130_fd_sc_hd__a21o_1 _17048_ (.A1(_09598_),
    .A2(_09599_),
    .B1(_09597_),
    .X(_09601_));
 sky130_fd_sc_hd__and3_1 _17049_ (.A(_09595_),
    .B(_09600_),
    .C(_09601_),
    .X(_09602_));
 sky130_fd_sc_hd__a21oi_1 _17050_ (.A1(_09600_),
    .A2(_09601_),
    .B1(_09595_),
    .Y(_09603_));
 sky130_fd_sc_hd__or3_1 _17051_ (.A(_09553_),
    .B(_09602_),
    .C(_09603_),
    .X(_09604_));
 sky130_fd_sc_hd__o21ai_1 _17052_ (.A1(_09602_),
    .A2(_09603_),
    .B1(_09553_),
    .Y(_09605_));
 sky130_fd_sc_hd__o21bai_1 _17053_ (.A1(_09553_),
    .A2(_09561_),
    .B1_N(net1117),
    .Y(_09606_));
 sky130_fd_sc_hd__nand3_1 _17054_ (.A(_09604_),
    .B(_09605_),
    .C(_09606_),
    .Y(_09607_));
 sky130_fd_sc_hd__a21o_1 _17055_ (.A1(_09604_),
    .A2(_09605_),
    .B1(_09606_),
    .X(_09608_));
 sky130_fd_sc_hd__and3_1 _17056_ (.A(_09594_),
    .B(_09607_),
    .C(_09608_),
    .X(_09609_));
 sky130_fd_sc_hd__a21oi_1 _17057_ (.A1(_09607_),
    .A2(_09608_),
    .B1(_09594_),
    .Y(_09610_));
 sky130_fd_sc_hd__or2_1 _17058_ (.A(_09609_),
    .B(_09610_),
    .X(_09611_));
 sky130_fd_sc_hd__a31o_1 _17059_ (.A1(_09562_),
    .A2(_09563_),
    .A3(_09564_),
    .B1(_09567_),
    .X(_09612_));
 sky130_fd_sc_hd__xnor2_2 _17060_ (.A(_09611_),
    .B(_09612_),
    .Y(_09613_));
 sky130_fd_sc_hd__xor2_1 _17061_ (.A(_09587_),
    .B(_09613_),
    .X(_09614_));
 sky130_fd_sc_hd__xnor2_1 _17062_ (.A(_09585_),
    .B(_09614_),
    .Y(_09615_));
 sky130_fd_sc_hd__or2_1 _17063_ (.A(_09584_),
    .B(_09615_),
    .X(_09616_));
 sky130_fd_sc_hd__nand2_1 _17064_ (.A(_09584_),
    .B(_09615_),
    .Y(_09617_));
 sky130_fd_sc_hd__nand2_1 _17065_ (.A(_09616_),
    .B(_09617_),
    .Y(_09618_));
 sky130_fd_sc_hd__xor2_1 _17066_ (.A(_09583_),
    .B(_09618_),
    .X(_09619_));
 sky130_fd_sc_hd__or2_1 _17067_ (.A(net1091),
    .B(_09494_),
    .X(_09620_));
 sky130_fd_sc_hd__o211a_1 _17068_ (.A1(_08870_),
    .A2(_09619_),
    .B1(_09620_),
    .C1(_09231_),
    .X(_00569_));
 sky130_fd_sc_hd__o21ai_1 _17069_ (.A1(_09583_),
    .A2(_09618_),
    .B1(_09616_),
    .Y(_09621_));
 sky130_fd_sc_hd__nand2_1 _17070_ (.A(_09585_),
    .B(_09614_),
    .Y(_09622_));
 sky130_fd_sc_hd__buf_4 _17071_ (.A(_09591_),
    .X(_09623_));
 sky130_fd_sc_hd__clkbuf_4 _17072_ (.A(_09623_),
    .X(_09624_));
 sky130_fd_sc_hd__clkbuf_4 _17073_ (.A(_09624_),
    .X(_09625_));
 sky130_fd_sc_hd__nor2_1 _17074_ (.A(_09625_),
    .B(_09592_),
    .Y(_09626_));
 sky130_fd_sc_hd__a21o_1 _17075_ (.A1(_09590_),
    .A2(_09593_),
    .B1(_09626_),
    .X(_09627_));
 sky130_fd_sc_hd__clkbuf_4 _17076_ (.A(_09459_),
    .X(_09628_));
 sky130_fd_sc_hd__clkbuf_4 _17077_ (.A(_09417_),
    .X(_09629_));
 sky130_fd_sc_hd__a21o_1 _17078_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[12] ),
    .A2(_09628_),
    .B1(_09629_),
    .X(_09630_));
 sky130_fd_sc_hd__clkbuf_8 _17079_ (.A(_09419_),
    .X(_09631_));
 sky130_fd_sc_hd__xnor2_2 _17080_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[13] ),
    .B(_09631_),
    .Y(_09632_));
 sky130_fd_sc_hd__xor2_2 _17081_ (.A(_09623_),
    .B(_09632_),
    .X(_09633_));
 sky130_fd_sc_hd__xor2_2 _17082_ (.A(_09630_),
    .B(_09633_),
    .X(_09634_));
 sky130_fd_sc_hd__a21bo_1 _17083_ (.A1(_09597_),
    .A2(_09599_),
    .B1_N(_09598_),
    .X(_09635_));
 sky130_fd_sc_hd__or4b_1 _17084_ (.A(_09361_),
    .B(_09377_),
    .C(_09215_),
    .D_N(net219),
    .X(_09636_));
 sky130_fd_sc_hd__a2bb2o_1 _17085_ (.A1_N(_09361_),
    .A2_N(_09215_),
    .B1(_09219_),
    .B2(_09213_),
    .X(_09637_));
 sky130_fd_sc_hd__nand3_1 _17086_ (.A(_09597_),
    .B(_09636_),
    .C(_09637_),
    .Y(_09638_));
 sky130_fd_sc_hd__a21o_1 _17087_ (.A1(_09636_),
    .A2(_09637_),
    .B1(_09597_),
    .X(_09639_));
 sky130_fd_sc_hd__and3_1 _17088_ (.A(_09635_),
    .B(_09638_),
    .C(_09639_),
    .X(_09640_));
 sky130_fd_sc_hd__a21oi_1 _17089_ (.A1(_09638_),
    .A2(_09639_),
    .B1(_09635_),
    .Y(_09641_));
 sky130_fd_sc_hd__or3_1 _17090_ (.A(_09553_),
    .B(_09640_),
    .C(_09641_),
    .X(_09642_));
 sky130_fd_sc_hd__o21ai_1 _17091_ (.A1(_09640_),
    .A2(_09641_),
    .B1(_09553_),
    .Y(_09643_));
 sky130_fd_sc_hd__o21bai_1 _17092_ (.A1(_09553_),
    .A2(_09603_),
    .B1_N(_09602_),
    .Y(_09644_));
 sky130_fd_sc_hd__nand3_1 _17093_ (.A(_09642_),
    .B(_09643_),
    .C(_09644_),
    .Y(_09645_));
 sky130_fd_sc_hd__a21o_1 _17094_ (.A1(_09642_),
    .A2(_09643_),
    .B1(_09644_),
    .X(_09646_));
 sky130_fd_sc_hd__nand3_1 _17095_ (.A(_09634_),
    .B(_09645_),
    .C(_09646_),
    .Y(_09647_));
 sky130_fd_sc_hd__a21o_1 _17096_ (.A1(_09645_),
    .A2(_09646_),
    .B1(_09634_),
    .X(_09648_));
 sky130_fd_sc_hd__a21bo_1 _17097_ (.A1(_09594_),
    .A2(_09608_),
    .B1_N(_09607_),
    .X(_09649_));
 sky130_fd_sc_hd__and3_1 _17098_ (.A(_09647_),
    .B(_09648_),
    .C(_09649_),
    .X(_09650_));
 sky130_fd_sc_hd__a21oi_1 _17099_ (.A1(_09647_),
    .A2(_09648_),
    .B1(_09649_),
    .Y(_09651_));
 sky130_fd_sc_hd__nor2_2 _17100_ (.A(_09650_),
    .B(_09651_),
    .Y(_09652_));
 sky130_fd_sc_hd__xnor2_2 _17101_ (.A(_09627_),
    .B(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__or2b_1 _17102_ (.A(_09611_),
    .B_N(_09612_),
    .X(_09654_));
 sky130_fd_sc_hd__nand2_1 _17103_ (.A(_09587_),
    .B(_09613_),
    .Y(_09655_));
 sky130_fd_sc_hd__nand2_1 _17104_ (.A(_09654_),
    .B(_09655_),
    .Y(_09656_));
 sky130_fd_sc_hd__xor2_1 _17105_ (.A(_09653_),
    .B(_09656_),
    .X(_09657_));
 sky130_fd_sc_hd__xnor2_1 _17106_ (.A(_09622_),
    .B(_09657_),
    .Y(_09658_));
 sky130_fd_sc_hd__nor2_1 _17107_ (.A(_09621_),
    .B(_09658_),
    .Y(_09659_));
 sky130_fd_sc_hd__a21o_1 _17108_ (.A1(_09621_),
    .A2(_09658_),
    .B1(_09292_),
    .X(_09660_));
 sky130_fd_sc_hd__o221a_1 _17109_ (.A1(net1049),
    .A2(_09266_),
    .B1(_09659_),
    .B2(_09660_),
    .C1(_07708_),
    .X(_00570_));
 sky130_fd_sc_hd__buf_4 _17110_ (.A(_04873_),
    .X(_09661_));
 sky130_fd_sc_hd__or2_1 _17111_ (.A(_09618_),
    .B(_09658_),
    .X(_09662_));
 sky130_fd_sc_hd__a21o_1 _17112_ (.A1(_09622_),
    .A2(_09616_),
    .B1(_09657_),
    .X(_09663_));
 sky130_fd_sc_hd__o21a_1 _17113_ (.A1(_09583_),
    .A2(_09662_),
    .B1(_09663_),
    .X(_09664_));
 sky130_fd_sc_hd__a21o_1 _17114_ (.A1(_09654_),
    .A2(_09655_),
    .B1(_09653_),
    .X(_09665_));
 sky130_fd_sc_hd__a21o_1 _17115_ (.A1(_09627_),
    .A2(_09652_),
    .B1(_09650_),
    .X(_09666_));
 sky130_fd_sc_hd__a21o_1 _17116_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[13] ),
    .A2(_09459_),
    .B1(_09417_),
    .X(_09667_));
 sky130_fd_sc_hd__xnor2_1 _17117_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[14] ),
    .B(_09419_),
    .Y(_09668_));
 sky130_fd_sc_hd__xor2_1 _17118_ (.A(_09623_),
    .B(_09668_),
    .X(_09669_));
 sky130_fd_sc_hd__xor2_1 _17119_ (.A(_09667_),
    .B(_09669_),
    .X(_09670_));
 sky130_fd_sc_hd__o21ba_1 _17120_ (.A1(_09553_),
    .A2(_09641_),
    .B1_N(_09640_),
    .X(_09671_));
 sky130_fd_sc_hd__nor2_1 _17121_ (.A(_09361_),
    .B(_09219_),
    .Y(_09672_));
 sky130_fd_sc_hd__a211o_1 _17122_ (.A1(_09213_),
    .A2(_09219_),
    .B1(_09597_),
    .C1(_09672_),
    .X(_09673_));
 sky130_fd_sc_hd__a21boi_1 _17123_ (.A1(_09597_),
    .A2(_09637_),
    .B1_N(_09636_),
    .Y(_09674_));
 sky130_fd_sc_hd__and3_1 _17124_ (.A(_09213_),
    .B(_09211_),
    .C(_09219_),
    .X(_09675_));
 sky130_fd_sc_hd__o211a_1 _17125_ (.A1(_09674_),
    .A2(_09675_),
    .B1(_09551_),
    .C1(_09552_),
    .X(_09676_));
 sky130_fd_sc_hd__a211oi_2 _17126_ (.A1(_09551_),
    .A2(_09552_),
    .B1(_09674_),
    .C1(_09675_),
    .Y(_09677_));
 sky130_fd_sc_hd__a21oi_2 _17127_ (.A1(_09551_),
    .A2(_09552_),
    .B1(_09673_),
    .Y(_09678_));
 sky130_fd_sc_hd__a211o_1 _17128_ (.A1(_09673_),
    .A2(_09676_),
    .B1(_09677_),
    .C1(_09678_),
    .X(_09679_));
 sky130_fd_sc_hd__xor2_1 _17129_ (.A(_09671_),
    .B(_09679_),
    .X(_09680_));
 sky130_fd_sc_hd__xnor2_1 _17130_ (.A(_09670_),
    .B(_09680_),
    .Y(_09681_));
 sky130_fd_sc_hd__a21boi_1 _17131_ (.A1(_09634_),
    .A2(_09646_),
    .B1_N(_09645_),
    .Y(_09682_));
 sky130_fd_sc_hd__xnor2_1 _17132_ (.A(_09681_),
    .B(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__nor2_1 _17133_ (.A(_09625_),
    .B(_09632_),
    .Y(_09684_));
 sky130_fd_sc_hd__a21o_1 _17134_ (.A1(_09630_),
    .A2(_09633_),
    .B1(_09684_),
    .X(_09685_));
 sky130_fd_sc_hd__or2b_1 _17135_ (.A(_09683_),
    .B_N(_09685_),
    .X(_09686_));
 sky130_fd_sc_hd__or2b_1 _17136_ (.A(_09685_),
    .B_N(_09683_),
    .X(_09687_));
 sky130_fd_sc_hd__nand2_1 _17137_ (.A(_09686_),
    .B(_09687_),
    .Y(_09688_));
 sky130_fd_sc_hd__xor2_1 _17138_ (.A(_09666_),
    .B(_09688_),
    .X(_09689_));
 sky130_fd_sc_hd__xor2_1 _17139_ (.A(_09665_),
    .B(_09689_),
    .X(_09690_));
 sky130_fd_sc_hd__and2b_1 _17140_ (.A_N(_09664_),
    .B(_09690_),
    .X(_09691_));
 sky130_fd_sc_hd__or2b_1 _17141_ (.A(_09690_),
    .B_N(_09664_),
    .X(_09692_));
 sky130_fd_sc_hd__nand2_1 _17142_ (.A(_06140_),
    .B(_09692_),
    .Y(_09693_));
 sky130_fd_sc_hd__a2bb2o_1 _17143_ (.A1_N(_09691_),
    .A2_N(_09693_),
    .B1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[14] ),
    .B2(_07816_),
    .X(_09694_));
 sky130_fd_sc_hd__and2_1 _17144_ (.A(_09661_),
    .B(_09694_),
    .X(_09695_));
 sky130_fd_sc_hd__clkbuf_1 _17145_ (.A(_09695_),
    .X(_00571_));
 sky130_fd_sc_hd__nor2_1 _17146_ (.A(_09665_),
    .B(_09689_),
    .Y(_09696_));
 sky130_fd_sc_hd__nor2_1 _17147_ (.A(_09696_),
    .B(_09691_),
    .Y(_09697_));
 sky130_fd_sc_hd__and2b_1 _17148_ (.A_N(_09688_),
    .B(_09666_),
    .X(_09698_));
 sky130_fd_sc_hd__or2_1 _17149_ (.A(_09681_),
    .B(_09682_),
    .X(_09699_));
 sky130_fd_sc_hd__nor2_1 _17150_ (.A(_09625_),
    .B(_09668_),
    .Y(_09700_));
 sky130_fd_sc_hd__a21o_1 _17151_ (.A1(_09667_),
    .A2(_09669_),
    .B1(_09700_),
    .X(_09701_));
 sky130_fd_sc_hd__nor2_1 _17152_ (.A(_09678_),
    .B(_09677_),
    .Y(_09702_));
 sky130_fd_sc_hd__a21o_1 _17153_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[14] ),
    .A2(_09459_),
    .B1(_09417_),
    .X(_09703_));
 sky130_fd_sc_hd__xnor2_1 _17154_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[15] ),
    .B(_09631_),
    .Y(_09704_));
 sky130_fd_sc_hd__xor2_1 _17155_ (.A(_09623_),
    .B(_09704_),
    .X(_09705_));
 sky130_fd_sc_hd__xnor2_1 _17156_ (.A(_09703_),
    .B(_09705_),
    .Y(_09706_));
 sky130_fd_sc_hd__xnor2_1 _17157_ (.A(_09702_),
    .B(_09706_),
    .Y(_09707_));
 sky130_fd_sc_hd__nor2_1 _17158_ (.A(_09671_),
    .B(_09679_),
    .Y(_09708_));
 sky130_fd_sc_hd__a21o_1 _17159_ (.A1(_09670_),
    .A2(_09680_),
    .B1(_09708_),
    .X(_09709_));
 sky130_fd_sc_hd__xor2_1 _17160_ (.A(_09707_),
    .B(_09709_),
    .X(_09710_));
 sky130_fd_sc_hd__xnor2_1 _17161_ (.A(_09701_),
    .B(_09710_),
    .Y(_09711_));
 sky130_fd_sc_hd__a21oi_1 _17162_ (.A1(_09699_),
    .A2(_09686_),
    .B1(_09711_),
    .Y(_09712_));
 sky130_fd_sc_hd__and3_1 _17163_ (.A(_09699_),
    .B(_09686_),
    .C(_09711_),
    .X(_09713_));
 sky130_fd_sc_hd__nor2_1 _17164_ (.A(_09712_),
    .B(_09713_),
    .Y(_09714_));
 sky130_fd_sc_hd__xor2_1 _17165_ (.A(_09698_),
    .B(_09714_),
    .X(_09715_));
 sky130_fd_sc_hd__and2_1 _17166_ (.A(_09697_),
    .B(_09715_),
    .X(_09716_));
 sky130_fd_sc_hd__o21ai_1 _17167_ (.A1(_09697_),
    .A2(_09715_),
    .B1(_06178_),
    .Y(_09717_));
 sky130_fd_sc_hd__o221a_1 _17168_ (.A1(net1055),
    .A2(_09266_),
    .B1(_09716_),
    .B2(_09717_),
    .C1(_07708_),
    .X(_00572_));
 sky130_fd_sc_hd__nand2_1 _17169_ (.A(_09690_),
    .B(_09715_),
    .Y(_09718_));
 sky130_fd_sc_hd__or2_1 _17170_ (.A(_09663_),
    .B(_09718_),
    .X(_09719_));
 sky130_fd_sc_hd__o21ai_1 _17171_ (.A1(_09698_),
    .A2(_09696_),
    .B1(_09714_),
    .Y(_09720_));
 sky130_fd_sc_hd__o311a_4 _17172_ (.A1(_09583_),
    .A2(_09662_),
    .A3(_09718_),
    .B1(_09719_),
    .C1(_09720_),
    .X(_09721_));
 sky130_fd_sc_hd__and2_1 _17173_ (.A(_09707_),
    .B(_09709_),
    .X(_09722_));
 sky130_fd_sc_hd__a21o_1 _17174_ (.A1(_09701_),
    .A2(_09710_),
    .B1(_09722_),
    .X(_09723_));
 sky130_fd_sc_hd__nor2_1 _17175_ (.A(_09625_),
    .B(_09704_),
    .Y(_09724_));
 sky130_fd_sc_hd__a21o_1 _17176_ (.A1(_09703_),
    .A2(_09705_),
    .B1(_09724_),
    .X(_09725_));
 sky130_fd_sc_hd__buf_2 _17177_ (.A(_09678_),
    .X(_09726_));
 sky130_fd_sc_hd__o21ba_1 _17178_ (.A1(_09726_),
    .A2(_09706_),
    .B1_N(_09677_),
    .X(_09727_));
 sky130_fd_sc_hd__a21o_1 _17179_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[15] ),
    .A2(_09459_),
    .B1(_09417_),
    .X(_09728_));
 sky130_fd_sc_hd__or3b_1 _17180_ (.A(_09417_),
    .B(_09418_),
    .C_N(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[16] ),
    .X(_09729_));
 sky130_fd_sc_hd__a21o_1 _17181_ (.A1(_09588_),
    .A2(_09459_),
    .B1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[16] ),
    .X(_09730_));
 sky130_fd_sc_hd__nand3b_1 _17182_ (.A_N(_09623_),
    .B(_09729_),
    .C(_09730_),
    .Y(_09731_));
 sky130_fd_sc_hd__a21bo_1 _17183_ (.A1(_09729_),
    .A2(_09730_),
    .B1_N(_09623_),
    .X(_09732_));
 sky130_fd_sc_hd__nand3_1 _17184_ (.A(_09728_),
    .B(_09731_),
    .C(_09732_),
    .Y(_09733_));
 sky130_fd_sc_hd__a21o_1 _17185_ (.A1(_09731_),
    .A2(_09732_),
    .B1(_09728_),
    .X(_09734_));
 sky130_fd_sc_hd__a21oi_1 _17186_ (.A1(_09733_),
    .A2(_09734_),
    .B1(_09726_),
    .Y(_09735_));
 sky130_fd_sc_hd__and3_1 _17187_ (.A(_09678_),
    .B(_09733_),
    .C(_09734_),
    .X(_09736_));
 sky130_fd_sc_hd__nor2_1 _17188_ (.A(_09735_),
    .B(_09736_),
    .Y(_09737_));
 sky130_fd_sc_hd__xnor2_1 _17189_ (.A(_09727_),
    .B(_09737_),
    .Y(_09738_));
 sky130_fd_sc_hd__xor2_1 _17190_ (.A(_09725_),
    .B(_09738_),
    .X(_09739_));
 sky130_fd_sc_hd__xnor2_1 _17191_ (.A(_09723_),
    .B(_09739_),
    .Y(_09740_));
 sky130_fd_sc_hd__nand2_1 _17192_ (.A(_09712_),
    .B(_09740_),
    .Y(_09741_));
 sky130_fd_sc_hd__or2_1 _17193_ (.A(_09712_),
    .B(_09740_),
    .X(_09742_));
 sky130_fd_sc_hd__nand2_1 _17194_ (.A(_09741_),
    .B(_09742_),
    .Y(_09743_));
 sky130_fd_sc_hd__or2_1 _17195_ (.A(_09721_),
    .B(_09743_),
    .X(_09744_));
 sky130_fd_sc_hd__nand2_1 _17196_ (.A(_09721_),
    .B(_09743_),
    .Y(_09745_));
 sky130_fd_sc_hd__and2_1 _17197_ (.A(_09744_),
    .B(_09745_),
    .X(_09746_));
 sky130_fd_sc_hd__or2_1 _17198_ (.A(net1080),
    .B(_09494_),
    .X(_09747_));
 sky130_fd_sc_hd__o211a_1 _17199_ (.A1(_08870_),
    .A2(_09746_),
    .B1(_09747_),
    .C1(_09231_),
    .X(_00573_));
 sky130_fd_sc_hd__or2b_1 _17200_ (.A(_09739_),
    .B_N(_09723_),
    .X(_09748_));
 sky130_fd_sc_hd__or2_1 _17201_ (.A(_09727_),
    .B(_09737_),
    .X(_09749_));
 sky130_fd_sc_hd__or2b_1 _17202_ (.A(_09738_),
    .B_N(_09725_),
    .X(_09750_));
 sky130_fd_sc_hd__nand2_1 _17203_ (.A(_09731_),
    .B(_09733_),
    .Y(_09751_));
 sky130_fd_sc_hd__and2_1 _17204_ (.A(_09588_),
    .B(_09729_),
    .X(_09752_));
 sky130_fd_sc_hd__or3b_1 _17205_ (.A(_09417_),
    .B(_09418_),
    .C_N(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[17] ),
    .X(_09753_));
 sky130_fd_sc_hd__a21o_1 _17206_ (.A1(_09588_),
    .A2(_09459_),
    .B1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[17] ),
    .X(_09754_));
 sky130_fd_sc_hd__nand3b_1 _17207_ (.A_N(_09623_),
    .B(_09753_),
    .C(_09754_),
    .Y(_09755_));
 sky130_fd_sc_hd__a21bo_1 _17208_ (.A1(_09753_),
    .A2(_09754_),
    .B1_N(_09623_),
    .X(_09756_));
 sky130_fd_sc_hd__nand2_1 _17209_ (.A(_09755_),
    .B(_09756_),
    .Y(_09757_));
 sky130_fd_sc_hd__xor2_2 _17210_ (.A(_09752_),
    .B(_09757_),
    .X(_09758_));
 sky130_fd_sc_hd__xnor2_1 _17211_ (.A(_09735_),
    .B(_09758_),
    .Y(_09759_));
 sky130_fd_sc_hd__xor2_1 _17212_ (.A(_09751_),
    .B(_09759_),
    .X(_09760_));
 sky130_fd_sc_hd__a21oi_1 _17213_ (.A1(_09749_),
    .A2(_09750_),
    .B1(_09760_),
    .Y(_09761_));
 sky130_fd_sc_hd__and3_1 _17214_ (.A(_09749_),
    .B(_09750_),
    .C(_09760_),
    .X(_09762_));
 sky130_fd_sc_hd__or2_1 _17215_ (.A(_09761_),
    .B(_09762_),
    .X(_09763_));
 sky130_fd_sc_hd__xor2_1 _17216_ (.A(_09748_),
    .B(_09763_),
    .X(_09764_));
 sky130_fd_sc_hd__a21oi_1 _17217_ (.A1(_09741_),
    .A2(_09744_),
    .B1(_09764_),
    .Y(_09765_));
 sky130_fd_sc_hd__a31o_1 _17218_ (.A1(_09741_),
    .A2(_09744_),
    .A3(_09764_),
    .B1(_07439_),
    .X(_09766_));
 sky130_fd_sc_hd__o221a_1 _17219_ (.A1(net1022),
    .A2(_09266_),
    .B1(_09765_),
    .B2(_09766_),
    .C1(_07708_),
    .X(_00574_));
 sky130_fd_sc_hd__a21oi_1 _17220_ (.A1(_09748_),
    .A2(_09741_),
    .B1(_09763_),
    .Y(_09767_));
 sky130_fd_sc_hd__or2b_1 _17221_ (.A(_09743_),
    .B_N(_09764_),
    .X(_09768_));
 sky130_fd_sc_hd__nor2_1 _17222_ (.A(net199),
    .B(_09768_),
    .Y(_09769_));
 sky130_fd_sc_hd__o21ai_1 _17223_ (.A1(_09752_),
    .A2(_09757_),
    .B1(_09755_),
    .Y(_09770_));
 sky130_fd_sc_hd__and2_1 _17224_ (.A(_09588_),
    .B(_09753_),
    .X(_09771_));
 sky130_fd_sc_hd__xnor2_2 _17225_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[18] ),
    .B(_09631_),
    .Y(_09772_));
 sky130_fd_sc_hd__xor2_2 _17226_ (.A(_09624_),
    .B(_09772_),
    .X(_09773_));
 sky130_fd_sc_hd__xnor2_2 _17227_ (.A(_09771_),
    .B(_09773_),
    .Y(_09774_));
 sky130_fd_sc_hd__or2_1 _17228_ (.A(_09726_),
    .B(_09758_),
    .X(_09775_));
 sky130_fd_sc_hd__xnor2_1 _17229_ (.A(_09774_),
    .B(_09775_),
    .Y(_09776_));
 sky130_fd_sc_hd__xnor2_1 _17230_ (.A(_09770_),
    .B(_09776_),
    .Y(_09777_));
 sky130_fd_sc_hd__nand2_1 _17231_ (.A(_09733_),
    .B(_09734_),
    .Y(_09778_));
 sky130_fd_sc_hd__or2b_1 _17232_ (.A(_09759_),
    .B_N(_09751_),
    .X(_09779_));
 sky130_fd_sc_hd__o21ai_1 _17233_ (.A1(_09778_),
    .A2(_09775_),
    .B1(_09779_),
    .Y(_09780_));
 sky130_fd_sc_hd__xnor2_1 _17234_ (.A(_09777_),
    .B(_09780_),
    .Y(_09781_));
 sky130_fd_sc_hd__xor2_1 _17235_ (.A(_09761_),
    .B(_09781_),
    .X(_09782_));
 sky130_fd_sc_hd__o21ai_1 _17236_ (.A1(_09767_),
    .A2(_09769_),
    .B1(_09782_),
    .Y(_09783_));
 sky130_fd_sc_hd__o31a_1 _17237_ (.A1(_09782_),
    .A2(_09767_),
    .A3(_09769_),
    .B1(_05311_),
    .X(_09784_));
 sky130_fd_sc_hd__a22o_1 _17238_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[18] ),
    .A2(_09496_),
    .B1(_09783_),
    .B2(_09784_),
    .X(_09785_));
 sky130_fd_sc_hd__and2_1 _17239_ (.A(_09661_),
    .B(_09785_),
    .X(_09786_));
 sky130_fd_sc_hd__clkbuf_1 _17240_ (.A(_09786_),
    .X(_00575_));
 sky130_fd_sc_hd__buf_6 _17241_ (.A(_05406_),
    .X(_09787_));
 sky130_fd_sc_hd__nand2_1 _17242_ (.A(_09761_),
    .B(_09781_),
    .Y(_09788_));
 sky130_fd_sc_hd__or2b_1 _17243_ (.A(_09777_),
    .B_N(_09780_),
    .X(_09789_));
 sky130_fd_sc_hd__or2b_1 _17244_ (.A(_09771_),
    .B_N(_09773_),
    .X(_09790_));
 sky130_fd_sc_hd__o21ai_1 _17245_ (.A1(_09625_),
    .A2(_09772_),
    .B1(_09790_),
    .Y(_09791_));
 sky130_fd_sc_hd__a21o_1 _17246_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[18] ),
    .A2(_09628_),
    .B1(_09629_),
    .X(_09792_));
 sky130_fd_sc_hd__xnor2_2 _17247_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[19] ),
    .B(_09631_),
    .Y(_09793_));
 sky130_fd_sc_hd__xor2_2 _17248_ (.A(_09623_),
    .B(_09793_),
    .X(_09794_));
 sky130_fd_sc_hd__xor2_2 _17249_ (.A(_09792_),
    .B(_09794_),
    .X(_09795_));
 sky130_fd_sc_hd__nor2_1 _17250_ (.A(_09726_),
    .B(_09774_),
    .Y(_09796_));
 sky130_fd_sc_hd__xor2_1 _17251_ (.A(_09795_),
    .B(_09796_),
    .X(_09797_));
 sky130_fd_sc_hd__xnor2_1 _17252_ (.A(_09791_),
    .B(_09797_),
    .Y(_09798_));
 sky130_fd_sc_hd__a22o_1 _17253_ (.A1(_09770_),
    .A2(_09776_),
    .B1(_09796_),
    .B2(_09758_),
    .X(_09799_));
 sky130_fd_sc_hd__xnor2_1 _17254_ (.A(_09798_),
    .B(_09799_),
    .Y(_09800_));
 sky130_fd_sc_hd__xnor2_1 _17255_ (.A(_09789_),
    .B(_09800_),
    .Y(_09801_));
 sky130_fd_sc_hd__a21oi_1 _17256_ (.A1(_09788_),
    .A2(_09783_),
    .B1(_09801_),
    .Y(_09802_));
 sky130_fd_sc_hd__and3_1 _17257_ (.A(_09788_),
    .B(_09783_),
    .C(_09801_),
    .X(_09803_));
 sky130_fd_sc_hd__buf_4 _17258_ (.A(_06701_),
    .X(_09804_));
 sky130_fd_sc_hd__or2_1 _17259_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[19] ),
    .B(_09804_),
    .X(_09805_));
 sky130_fd_sc_hd__clkbuf_8 _17260_ (.A(_04869_),
    .X(_09806_));
 sky130_fd_sc_hd__o311a_1 _17261_ (.A1(_09787_),
    .A2(_09802_),
    .A3(_09803_),
    .B1(_09805_),
    .C1(_09806_),
    .X(_00576_));
 sky130_fd_sc_hd__and2b_1 _17262_ (.A_N(_09798_),
    .B(_09799_),
    .X(_09807_));
 sky130_fd_sc_hd__nand2_1 _17263_ (.A(_09791_),
    .B(_09797_),
    .Y(_09808_));
 sky130_fd_sc_hd__nor2_1 _17264_ (.A(_09726_),
    .B(_09795_),
    .Y(_09809_));
 sky130_fd_sc_hd__nand2_1 _17265_ (.A(_09774_),
    .B(_09809_),
    .Y(_09810_));
 sky130_fd_sc_hd__nor2_1 _17266_ (.A(_09625_),
    .B(_09793_),
    .Y(_09811_));
 sky130_fd_sc_hd__a21o_1 _17267_ (.A1(_09792_),
    .A2(_09794_),
    .B1(_09811_),
    .X(_09812_));
 sky130_fd_sc_hd__a21o_1 _17268_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[19] ),
    .A2(_09628_),
    .B1(_09629_),
    .X(_09813_));
 sky130_fd_sc_hd__xnor2_2 _17269_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[20] ),
    .B(_09631_),
    .Y(_09814_));
 sky130_fd_sc_hd__xor2_2 _17270_ (.A(_09624_),
    .B(_09814_),
    .X(_09815_));
 sky130_fd_sc_hd__xor2_2 _17271_ (.A(_09813_),
    .B(_09815_),
    .X(_09816_));
 sky130_fd_sc_hd__xor2_1 _17272_ (.A(_09816_),
    .B(_09809_),
    .X(_09817_));
 sky130_fd_sc_hd__xnor2_1 _17273_ (.A(_09812_),
    .B(_09817_),
    .Y(_09818_));
 sky130_fd_sc_hd__a21o_1 _17274_ (.A1(_09808_),
    .A2(_09810_),
    .B1(_09818_),
    .X(_09819_));
 sky130_fd_sc_hd__nand3_1 _17275_ (.A(_09808_),
    .B(_09818_),
    .C(_09810_),
    .Y(_09820_));
 sky130_fd_sc_hd__and2_1 _17276_ (.A(_09819_),
    .B(_09820_),
    .X(_09821_));
 sky130_fd_sc_hd__xnor2_1 _17277_ (.A(_09807_),
    .B(_09821_),
    .Y(_09822_));
 sky130_fd_sc_hd__and2_1 _17278_ (.A(_09782_),
    .B(_09801_),
    .X(_09823_));
 sky130_fd_sc_hd__or2b_2 _17279_ (.A(_09768_),
    .B_N(_09823_),
    .X(_09824_));
 sky130_fd_sc_hd__nand2_1 _17280_ (.A(_09789_),
    .B(_09788_),
    .Y(_09825_));
 sky130_fd_sc_hd__a22o_1 _17281_ (.A1(_09767_),
    .A2(_09823_),
    .B1(_09825_),
    .B2(_09800_),
    .X(_09826_));
 sky130_fd_sc_hd__o21bai_2 _17282_ (.A1(_09721_),
    .A2(_09824_),
    .B1_N(_09826_),
    .Y(_09827_));
 sky130_fd_sc_hd__xnor2_1 _17283_ (.A(_09822_),
    .B(_09827_),
    .Y(_09828_));
 sky130_fd_sc_hd__or2_1 _17284_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[20] ),
    .B(_09494_),
    .X(_09829_));
 sky130_fd_sc_hd__o211a_1 _17285_ (.A1(_08870_),
    .A2(_09828_),
    .B1(_09829_),
    .C1(_09231_),
    .X(_00577_));
 sky130_fd_sc_hd__nand2_1 _17286_ (.A(_09807_),
    .B(_09821_),
    .Y(_09830_));
 sky130_fd_sc_hd__or2b_1 _17287_ (.A(_09822_),
    .B_N(_09827_),
    .X(_09831_));
 sky130_fd_sc_hd__nor2_1 _17288_ (.A(_09625_),
    .B(_09814_),
    .Y(_09832_));
 sky130_fd_sc_hd__a21o_1 _17289_ (.A1(_09813_),
    .A2(_09815_),
    .B1(_09832_),
    .X(_09833_));
 sky130_fd_sc_hd__a21o_1 _17290_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[20] ),
    .A2(_09628_),
    .B1(_09629_),
    .X(_09834_));
 sky130_fd_sc_hd__xnor2_1 _17291_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[21] ),
    .B(_09631_),
    .Y(_09835_));
 sky130_fd_sc_hd__or2_1 _17292_ (.A(_09623_),
    .B(_09835_),
    .X(_09836_));
 sky130_fd_sc_hd__nand2_1 _17293_ (.A(_09624_),
    .B(_09835_),
    .Y(_09837_));
 sky130_fd_sc_hd__and2_2 _17294_ (.A(_09836_),
    .B(_09837_),
    .X(_09838_));
 sky130_fd_sc_hd__xor2_2 _17295_ (.A(_09834_),
    .B(_09838_),
    .X(_09839_));
 sky130_fd_sc_hd__nor2_1 _17296_ (.A(_09726_),
    .B(_09816_),
    .Y(_09840_));
 sky130_fd_sc_hd__xor2_1 _17297_ (.A(_09839_),
    .B(_09840_),
    .X(_09841_));
 sky130_fd_sc_hd__xnor2_1 _17298_ (.A(_09833_),
    .B(_09841_),
    .Y(_09842_));
 sky130_fd_sc_hd__a22oi_1 _17299_ (.A1(_09812_),
    .A2(_09817_),
    .B1(_09840_),
    .B2(_09795_),
    .Y(_09843_));
 sky130_fd_sc_hd__nor2_1 _17300_ (.A(_09842_),
    .B(_09843_),
    .Y(_09844_));
 sky130_fd_sc_hd__and2_1 _17301_ (.A(_09842_),
    .B(_09843_),
    .X(_09845_));
 sky130_fd_sc_hd__nor2_1 _17302_ (.A(_09844_),
    .B(_09845_),
    .Y(_09846_));
 sky130_fd_sc_hd__xnor2_1 _17303_ (.A(_09819_),
    .B(_09846_),
    .Y(_09847_));
 sky130_fd_sc_hd__a21oi_1 _17304_ (.A1(_09830_),
    .A2(_09831_),
    .B1(_09847_),
    .Y(_09848_));
 sky130_fd_sc_hd__a31o_1 _17305_ (.A1(_09830_),
    .A2(_09831_),
    .A3(_09847_),
    .B1(_07439_),
    .X(_09849_));
 sky130_fd_sc_hd__o221a_1 _17306_ (.A1(net1050),
    .A2(_09266_),
    .B1(_09848_),
    .B2(_09849_),
    .C1(_07708_),
    .X(_00578_));
 sky130_fd_sc_hd__and2b_1 _17307_ (.A_N(_09822_),
    .B(_09847_),
    .X(_09850_));
 sky130_fd_sc_hd__a21boi_1 _17308_ (.A1(_09819_),
    .A2(_09830_),
    .B1_N(_09846_),
    .Y(_09851_));
 sky130_fd_sc_hd__a21oi_1 _17309_ (.A1(_09827_),
    .A2(_09850_),
    .B1(_09851_),
    .Y(_09852_));
 sky130_fd_sc_hd__a21bo_1 _17310_ (.A1(_09834_),
    .A2(_09837_),
    .B1_N(_09836_),
    .X(_09853_));
 sky130_fd_sc_hd__a21oi_2 _17311_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[21] ),
    .A2(_09628_),
    .B1(_09629_),
    .Y(_09854_));
 sky130_fd_sc_hd__xnor2_2 _17312_ (.A(_09838_),
    .B(_09854_),
    .Y(_09855_));
 sky130_fd_sc_hd__nor2_1 _17313_ (.A(_09726_),
    .B(_09839_),
    .Y(_09856_));
 sky130_fd_sc_hd__xor2_1 _17314_ (.A(_09855_),
    .B(_09856_),
    .X(_09857_));
 sky130_fd_sc_hd__xnor2_1 _17315_ (.A(_09853_),
    .B(_09857_),
    .Y(_09858_));
 sky130_fd_sc_hd__a22o_1 _17316_ (.A1(_09833_),
    .A2(_09841_),
    .B1(_09856_),
    .B2(_09816_),
    .X(_09859_));
 sky130_fd_sc_hd__xnor2_1 _17317_ (.A(_09858_),
    .B(_09859_),
    .Y(_09860_));
 sky130_fd_sc_hd__or2_1 _17318_ (.A(_09844_),
    .B(_09860_),
    .X(_09861_));
 sky130_fd_sc_hd__nand2_1 _17319_ (.A(_09844_),
    .B(_09860_),
    .Y(_09862_));
 sky130_fd_sc_hd__nand2_1 _17320_ (.A(_09861_),
    .B(_09862_),
    .Y(_09863_));
 sky130_fd_sc_hd__nor2_1 _17321_ (.A(_05399_),
    .B(_09863_),
    .Y(_09864_));
 sky130_fd_sc_hd__a22o_1 _17322_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[22] ),
    .A2(_09496_),
    .B1(_09852_),
    .B2(_09864_),
    .X(_09865_));
 sky130_fd_sc_hd__and2_1 _17323_ (.A(_09661_),
    .B(_09865_),
    .X(_09866_));
 sky130_fd_sc_hd__clkbuf_1 _17324_ (.A(_09866_),
    .X(_00579_));
 sky130_fd_sc_hd__or2b_1 _17325_ (.A(_09858_),
    .B_N(_09859_),
    .X(_09867_));
 sky130_fd_sc_hd__nand2_1 _17326_ (.A(_09853_),
    .B(_09857_),
    .Y(_09868_));
 sky130_fd_sc_hd__nor2_1 _17327_ (.A(_09726_),
    .B(_09855_),
    .Y(_09869_));
 sky130_fd_sc_hd__nand2_1 _17328_ (.A(_09839_),
    .B(_09869_),
    .Y(_09870_));
 sky130_fd_sc_hd__a21o_1 _17329_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[21] ),
    .A2(_09628_),
    .B1(_09629_),
    .X(_09871_));
 sky130_fd_sc_hd__a21bo_1 _17330_ (.A1(_09837_),
    .A2(_09871_),
    .B1_N(_09836_),
    .X(_09872_));
 sky130_fd_sc_hd__xnor2_1 _17331_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[23] ),
    .B(_09631_),
    .Y(_09873_));
 sky130_fd_sc_hd__nor2_1 _17332_ (.A(_09624_),
    .B(_09873_),
    .Y(_09874_));
 sky130_fd_sc_hd__nand2_1 _17333_ (.A(_09624_),
    .B(_09873_),
    .Y(_09875_));
 sky130_fd_sc_hd__and2b_1 _17334_ (.A_N(_09874_),
    .B(_09875_),
    .X(_09876_));
 sky130_fd_sc_hd__xnor2_2 _17335_ (.A(_09854_),
    .B(_09876_),
    .Y(_09877_));
 sky130_fd_sc_hd__xor2_1 _17336_ (.A(_09877_),
    .B(_09869_),
    .X(_09878_));
 sky130_fd_sc_hd__xnor2_1 _17337_ (.A(_09872_),
    .B(_09878_),
    .Y(_09879_));
 sky130_fd_sc_hd__a21o_1 _17338_ (.A1(_09868_),
    .A2(_09870_),
    .B1(_09879_),
    .X(_09880_));
 sky130_fd_sc_hd__nand3_1 _17339_ (.A(_09868_),
    .B(_09879_),
    .C(_09870_),
    .Y(_09881_));
 sky130_fd_sc_hd__and2_1 _17340_ (.A(_09880_),
    .B(_09881_),
    .X(_09882_));
 sky130_fd_sc_hd__xnor2_1 _17341_ (.A(_09867_),
    .B(_09882_),
    .Y(_09883_));
 sky130_fd_sc_hd__a21oi_1 _17342_ (.A1(_09852_),
    .A2(_09862_),
    .B1(_09883_),
    .Y(_09884_));
 sky130_fd_sc_hd__a31o_1 _17343_ (.A1(_09852_),
    .A2(_09862_),
    .A3(_09883_),
    .B1(_07439_),
    .X(_09885_));
 sky130_fd_sc_hd__clkbuf_8 _17344_ (.A(_07707_),
    .X(_09886_));
 sky130_fd_sc_hd__o221a_1 _17345_ (.A1(net1047),
    .A2(_09266_),
    .B1(_09884_),
    .B2(_09885_),
    .C1(_09886_),
    .X(_00580_));
 sky130_fd_sc_hd__and2b_1 _17346_ (.A_N(_09863_),
    .B(_09883_),
    .X(_09887_));
 sky130_fd_sc_hd__nand2_1 _17347_ (.A(_09850_),
    .B(_09887_),
    .Y(_09888_));
 sky130_fd_sc_hd__nand2_1 _17348_ (.A(_09867_),
    .B(_09862_),
    .Y(_09889_));
 sky130_fd_sc_hd__a21o_1 _17349_ (.A1(_09826_),
    .A2(_09850_),
    .B1(_09851_),
    .X(_09890_));
 sky130_fd_sc_hd__a22oi_2 _17350_ (.A1(_09882_),
    .A2(_09889_),
    .B1(_09887_),
    .B2(_09890_),
    .Y(_09891_));
 sky130_fd_sc_hd__o31ai_4 _17351_ (.A1(_09721_),
    .A2(_09824_),
    .A3(_09888_),
    .B1(_09891_),
    .Y(_09892_));
 sky130_fd_sc_hd__a21o_1 _17352_ (.A1(_09871_),
    .A2(_09875_),
    .B1(_09874_),
    .X(_09893_));
 sky130_fd_sc_hd__a21o_1 _17353_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[23] ),
    .A2(_09628_),
    .B1(_09629_),
    .X(_09894_));
 sky130_fd_sc_hd__xnor2_1 _17354_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[24] ),
    .B(_09631_),
    .Y(_09895_));
 sky130_fd_sc_hd__nor2_1 _17355_ (.A(_09624_),
    .B(_09895_),
    .Y(_09896_));
 sky130_fd_sc_hd__nand2_1 _17356_ (.A(_09625_),
    .B(_09895_),
    .Y(_09897_));
 sky130_fd_sc_hd__and2b_1 _17357_ (.A_N(_09896_),
    .B(_09897_),
    .X(_09898_));
 sky130_fd_sc_hd__xor2_2 _17358_ (.A(_09894_),
    .B(_09898_),
    .X(_09899_));
 sky130_fd_sc_hd__nor2_1 _17359_ (.A(_09726_),
    .B(_09877_),
    .Y(_09900_));
 sky130_fd_sc_hd__xnor2_2 _17360_ (.A(_09899_),
    .B(_09900_),
    .Y(_09901_));
 sky130_fd_sc_hd__xnor2_2 _17361_ (.A(_09893_),
    .B(_09901_),
    .Y(_09902_));
 sky130_fd_sc_hd__a22o_1 _17362_ (.A1(_09872_),
    .A2(_09878_),
    .B1(_09900_),
    .B2(_09855_),
    .X(_09903_));
 sky130_fd_sc_hd__xor2_2 _17363_ (.A(_09902_),
    .B(_09903_),
    .X(_09904_));
 sky130_fd_sc_hd__xnor2_2 _17364_ (.A(_09880_),
    .B(_09904_),
    .Y(_09905_));
 sky130_fd_sc_hd__xor2_1 _17365_ (.A(net252),
    .B(_09905_),
    .X(_09906_));
 sky130_fd_sc_hd__or2_1 _17366_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[24] ),
    .B(_09494_),
    .X(_09907_));
 sky130_fd_sc_hd__o211a_1 _17367_ (.A1(_08870_),
    .A2(_09906_),
    .B1(_09907_),
    .C1(_09231_),
    .X(_00581_));
 sky130_fd_sc_hd__or2b_1 _17368_ (.A(_09880_),
    .B_N(_09904_),
    .X(_09908_));
 sky130_fd_sc_hd__nand2_1 _17369_ (.A(_09892_),
    .B(_09905_),
    .Y(_09909_));
 sky130_fd_sc_hd__nand2_1 _17370_ (.A(_09902_),
    .B(_09903_),
    .Y(_09910_));
 sky130_fd_sc_hd__a21o_1 _17371_ (.A1(_09894_),
    .A2(_09897_),
    .B1(_09896_),
    .X(_09911_));
 sky130_fd_sc_hd__xnor2_1 _17372_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[25] ),
    .B(_09631_),
    .Y(_09912_));
 sky130_fd_sc_hd__or2_2 _17373_ (.A(_09624_),
    .B(_09912_),
    .X(_09913_));
 sky130_fd_sc_hd__nand2_1 _17374_ (.A(_09624_),
    .B(_09912_),
    .Y(_09914_));
 sky130_fd_sc_hd__nand2_2 _17375_ (.A(_09913_),
    .B(_09914_),
    .Y(_09915_));
 sky130_fd_sc_hd__a21oi_1 _17376_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[24] ),
    .A2(_09628_),
    .B1(_09629_),
    .Y(_09916_));
 sky130_fd_sc_hd__xor2_1 _17377_ (.A(_09915_),
    .B(_09916_),
    .X(_09917_));
 sky130_fd_sc_hd__inv_2 _17378_ (.A(_09917_),
    .Y(_09918_));
 sky130_fd_sc_hd__buf_2 _17379_ (.A(_09726_),
    .X(_09919_));
 sky130_fd_sc_hd__nor2_1 _17380_ (.A(_09919_),
    .B(_09899_),
    .Y(_09920_));
 sky130_fd_sc_hd__xnor2_1 _17381_ (.A(_09918_),
    .B(_09920_),
    .Y(_09921_));
 sky130_fd_sc_hd__xnor2_1 _17382_ (.A(_09911_),
    .B(_09921_),
    .Y(_09922_));
 sky130_fd_sc_hd__and2b_1 _17383_ (.A_N(_09901_),
    .B(_09893_),
    .X(_09923_));
 sky130_fd_sc_hd__a21oi_1 _17384_ (.A1(_09877_),
    .A2(_09920_),
    .B1(_09923_),
    .Y(_09924_));
 sky130_fd_sc_hd__xor2_1 _17385_ (.A(_09922_),
    .B(_09924_),
    .X(_09925_));
 sky130_fd_sc_hd__xnor2_1 _17386_ (.A(_09910_),
    .B(_09925_),
    .Y(_09926_));
 sky130_fd_sc_hd__a21oi_1 _17387_ (.A1(_09908_),
    .A2(_09909_),
    .B1(_09926_),
    .Y(_09927_));
 sky130_fd_sc_hd__a31o_1 _17388_ (.A1(_09908_),
    .A2(_09909_),
    .A3(_09926_),
    .B1(_07439_),
    .X(_09928_));
 sky130_fd_sc_hd__o221a_1 _17389_ (.A1(net1051),
    .A2(_09266_),
    .B1(_09927_),
    .B2(_09928_),
    .C1(_09886_),
    .X(_00582_));
 sky130_fd_sc_hd__nand2_1 _17390_ (.A(_09905_),
    .B(_09926_),
    .Y(_09929_));
 sky130_fd_sc_hd__inv_2 _17391_ (.A(_09929_),
    .Y(_09930_));
 sky130_fd_sc_hd__a21boi_1 _17392_ (.A1(_09910_),
    .A2(_09908_),
    .B1_N(_09925_),
    .Y(_09931_));
 sky130_fd_sc_hd__a21oi_1 _17393_ (.A1(_09892_),
    .A2(_09930_),
    .B1(_09931_),
    .Y(_09932_));
 sky130_fd_sc_hd__nor2_1 _17394_ (.A(_09922_),
    .B(_09924_),
    .Y(_09933_));
 sky130_fd_sc_hd__or2_1 _17395_ (.A(_09915_),
    .B(_09916_),
    .X(_09934_));
 sky130_fd_sc_hd__a21oi_2 _17396_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[25] ),
    .A2(_09628_),
    .B1(_09629_),
    .Y(_09935_));
 sky130_fd_sc_hd__inv_2 _17397_ (.A(_09935_),
    .Y(_09936_));
 sky130_fd_sc_hd__xnor2_2 _17398_ (.A(_09915_),
    .B(_09936_),
    .Y(_09937_));
 sky130_fd_sc_hd__nor2_1 _17399_ (.A(_09919_),
    .B(_09917_),
    .Y(_09938_));
 sky130_fd_sc_hd__xnor2_1 _17400_ (.A(_09937_),
    .B(_09938_),
    .Y(_09939_));
 sky130_fd_sc_hd__a21o_1 _17401_ (.A1(_09913_),
    .A2(_09934_),
    .B1(_09939_),
    .X(_09940_));
 sky130_fd_sc_hd__nand3_1 _17402_ (.A(_09913_),
    .B(_09934_),
    .C(_09939_),
    .Y(_09941_));
 sky130_fd_sc_hd__nand2_1 _17403_ (.A(_09940_),
    .B(_09941_),
    .Y(_09942_));
 sky130_fd_sc_hd__a22o_1 _17404_ (.A1(_09911_),
    .A2(_09921_),
    .B1(_09938_),
    .B2(_09899_),
    .X(_09943_));
 sky130_fd_sc_hd__xnor2_1 _17405_ (.A(_09942_),
    .B(_09943_),
    .Y(_09944_));
 sky130_fd_sc_hd__or2_1 _17406_ (.A(_09933_),
    .B(_09944_),
    .X(_09945_));
 sky130_fd_sc_hd__nand2_1 _17407_ (.A(_09933_),
    .B(_09944_),
    .Y(_09946_));
 sky130_fd_sc_hd__nand2_1 _17408_ (.A(_09945_),
    .B(_09946_),
    .Y(_09947_));
 sky130_fd_sc_hd__nor2_1 _17409_ (.A(_05405_),
    .B(_09947_),
    .Y(_09948_));
 sky130_fd_sc_hd__a22o_1 _17410_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[26] ),
    .A2(_09496_),
    .B1(_09932_),
    .B2(_09948_),
    .X(_09949_));
 sky130_fd_sc_hd__and2_1 _17411_ (.A(_09661_),
    .B(_09949_),
    .X(_09950_));
 sky130_fd_sc_hd__clkbuf_1 _17412_ (.A(_09950_),
    .X(_00583_));
 sky130_fd_sc_hd__or2b_1 _17413_ (.A(_09942_),
    .B_N(_09943_),
    .X(_09951_));
 sky130_fd_sc_hd__o21a_1 _17414_ (.A1(_09915_),
    .A2(_09935_),
    .B1(_09913_),
    .X(_09952_));
 sky130_fd_sc_hd__xnor2_1 _17415_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[27] ),
    .B(_09631_),
    .Y(_09953_));
 sky130_fd_sc_hd__or2_1 _17416_ (.A(_09624_),
    .B(_09953_),
    .X(_09954_));
 sky130_fd_sc_hd__nand2_1 _17417_ (.A(_09625_),
    .B(_09953_),
    .Y(_09955_));
 sky130_fd_sc_hd__nand2_2 _17418_ (.A(_09954_),
    .B(_09955_),
    .Y(_09956_));
 sky130_fd_sc_hd__xnor2_2 _17419_ (.A(_09936_),
    .B(_09956_),
    .Y(_09957_));
 sky130_fd_sc_hd__nor2_1 _17420_ (.A(_09919_),
    .B(_09957_),
    .Y(_09958_));
 sky130_fd_sc_hd__and2_1 _17421_ (.A(_09919_),
    .B(_09957_),
    .X(_09959_));
 sky130_fd_sc_hd__nor2_1 _17422_ (.A(_09958_),
    .B(_09959_),
    .Y(_09960_));
 sky130_fd_sc_hd__xnor2_1 _17423_ (.A(_09935_),
    .B(_09956_),
    .Y(_09961_));
 sky130_fd_sc_hd__mux2_1 _17424_ (.A0(_09960_),
    .A1(_09961_),
    .S(_09937_),
    .X(_09962_));
 sky130_fd_sc_hd__xnor2_1 _17425_ (.A(_09952_),
    .B(_09962_),
    .Y(_09963_));
 sky130_fd_sc_hd__o31a_1 _17426_ (.A1(_09919_),
    .A2(_09918_),
    .A3(_09937_),
    .B1(_09940_),
    .X(_09964_));
 sky130_fd_sc_hd__nor2_1 _17427_ (.A(_09963_),
    .B(_09964_),
    .Y(_09965_));
 sky130_fd_sc_hd__and2_1 _17428_ (.A(_09963_),
    .B(_09964_),
    .X(_09966_));
 sky130_fd_sc_hd__nor2_1 _17429_ (.A(_09965_),
    .B(_09966_),
    .Y(_09967_));
 sky130_fd_sc_hd__xnor2_1 _17430_ (.A(_09951_),
    .B(_09967_),
    .Y(_09968_));
 sky130_fd_sc_hd__a21oi_1 _17431_ (.A1(_09932_),
    .A2(_09946_),
    .B1(_09968_),
    .Y(_09969_));
 sky130_fd_sc_hd__and3_1 _17432_ (.A(_09932_),
    .B(_09946_),
    .C(_09968_),
    .X(_09970_));
 sky130_fd_sc_hd__or2_1 _17433_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[27] ),
    .B(_05316_),
    .X(_09971_));
 sky130_fd_sc_hd__o311a_1 _17434_ (.A1(_09787_),
    .A2(_09969_),
    .A3(_09970_),
    .B1(_09971_),
    .C1(_09806_),
    .X(_00584_));
 sky130_fd_sc_hd__o21a_1 _17435_ (.A1(_09935_),
    .A2(_09956_),
    .B1(_09954_),
    .X(_09972_));
 sky130_fd_sc_hd__a21oi_1 _17436_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[27] ),
    .A2(_09628_),
    .B1(_09629_),
    .Y(_09973_));
 sky130_fd_sc_hd__or2_1 _17437_ (.A(_09915_),
    .B(_09973_),
    .X(_09974_));
 sky130_fd_sc_hd__nand2_1 _17438_ (.A(_09915_),
    .B(_09973_),
    .Y(_09975_));
 sky130_fd_sc_hd__nand2_1 _17439_ (.A(_09974_),
    .B(_09975_),
    .Y(_09976_));
 sky130_fd_sc_hd__xnor2_1 _17440_ (.A(_09958_),
    .B(_09976_),
    .Y(_09977_));
 sky130_fd_sc_hd__and2b_1 _17441_ (.A_N(_09972_),
    .B(_09977_),
    .X(_09978_));
 sky130_fd_sc_hd__and2b_1 _17442_ (.A_N(_09977_),
    .B(_09972_),
    .X(_09979_));
 sky130_fd_sc_hd__or2_1 _17443_ (.A(_09978_),
    .B(_09979_),
    .X(_09980_));
 sky130_fd_sc_hd__or3b_1 _17444_ (.A(_09919_),
    .B(_09957_),
    .C_N(_09937_),
    .X(_09981_));
 sky130_fd_sc_hd__o21ai_1 _17445_ (.A1(_09952_),
    .A2(_09962_),
    .B1(_09981_),
    .Y(_09982_));
 sky130_fd_sc_hd__xnor2_1 _17446_ (.A(_09980_),
    .B(_09982_),
    .Y(_09983_));
 sky130_fd_sc_hd__or2_1 _17447_ (.A(_09965_),
    .B(_09983_),
    .X(_09984_));
 sky130_fd_sc_hd__nand2_1 _17448_ (.A(_09965_),
    .B(_09983_),
    .Y(_09985_));
 sky130_fd_sc_hd__inv_2 _17449_ (.A(_09947_),
    .Y(_09986_));
 sky130_fd_sc_hd__and3_1 _17450_ (.A(_09930_),
    .B(_09986_),
    .C(_09968_),
    .X(_09987_));
 sky130_fd_sc_hd__nand2_1 _17451_ (.A(_09951_),
    .B(_09946_),
    .Y(_09988_));
 sky130_fd_sc_hd__a32o_1 _17452_ (.A1(_09931_),
    .A2(_09986_),
    .A3(_09968_),
    .B1(_09988_),
    .B2(_09967_),
    .X(_09989_));
 sky130_fd_sc_hd__a21oi_2 _17453_ (.A1(_09892_),
    .A2(_09987_),
    .B1(_09989_),
    .Y(_09990_));
 sky130_fd_sc_hd__a31o_1 _17454_ (.A1(_09984_),
    .A2(_09985_),
    .A3(_09990_),
    .B1(_05732_),
    .X(_09991_));
 sky130_fd_sc_hd__o211a_1 _17455_ (.A1(net1030),
    .A2(_08183_),
    .B1(_09991_),
    .C1(_09231_),
    .X(_00585_));
 sky130_fd_sc_hd__or2b_1 _17456_ (.A(_09980_),
    .B_N(_09982_),
    .X(_09992_));
 sky130_fd_sc_hd__and3b_1 _17457_ (.A_N(_09919_),
    .B(_09957_),
    .C(_09976_),
    .X(_09993_));
 sky130_fd_sc_hd__mux2_1 _17458_ (.A0(_09961_),
    .A1(_09960_),
    .S(_09976_),
    .X(_09994_));
 sky130_fd_sc_hd__a21o_1 _17459_ (.A1(_09913_),
    .A2(_09974_),
    .B1(_09994_),
    .X(_09995_));
 sky130_fd_sc_hd__nand3_1 _17460_ (.A(_09913_),
    .B(_09974_),
    .C(_09994_),
    .Y(_09996_));
 sky130_fd_sc_hd__and2_1 _17461_ (.A(_09995_),
    .B(_09996_),
    .X(_09997_));
 sky130_fd_sc_hd__o21a_1 _17462_ (.A1(_09978_),
    .A2(_09993_),
    .B1(_09997_),
    .X(_09998_));
 sky130_fd_sc_hd__nor3_1 _17463_ (.A(_09978_),
    .B(_09997_),
    .C(_09993_),
    .Y(_09999_));
 sky130_fd_sc_hd__a211o_1 _17464_ (.A1(_09992_),
    .A2(_09985_),
    .B1(_09998_),
    .C1(_09999_),
    .X(_10000_));
 sky130_fd_sc_hd__or3_1 _17465_ (.A(_09919_),
    .B(_09957_),
    .C(_09976_),
    .X(_10001_));
 sky130_fd_sc_hd__mux2_1 _17466_ (.A0(_09936_),
    .A1(_09956_),
    .S(_09919_),
    .X(_10002_));
 sky130_fd_sc_hd__xnor2_1 _17467_ (.A(_09972_),
    .B(_10002_),
    .Y(_10003_));
 sky130_fd_sc_hd__xnor2_1 _17468_ (.A(_09973_),
    .B(_10003_),
    .Y(_10004_));
 sky130_fd_sc_hd__a21o_1 _17469_ (.A1(_10001_),
    .A2(_09995_),
    .B1(_10004_),
    .X(_10005_));
 sky130_fd_sc_hd__nand3_1 _17470_ (.A(_10001_),
    .B(_09995_),
    .C(_10004_),
    .Y(_10006_));
 sky130_fd_sc_hd__and2_1 _17471_ (.A(_10005_),
    .B(_10006_),
    .X(_10007_));
 sky130_fd_sc_hd__nand2_1 _17472_ (.A(_09998_),
    .B(_10007_),
    .Y(_10008_));
 sky130_fd_sc_hd__or2_1 _17473_ (.A(_09998_),
    .B(_10007_),
    .X(_10009_));
 sky130_fd_sc_hd__and4_1 _17474_ (.A(_09990_),
    .B(_10000_),
    .C(_10008_),
    .D(_10009_),
    .X(_10010_));
 sky130_fd_sc_hd__or2_1 _17475_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[29] ),
    .B(_09494_),
    .X(_10011_));
 sky130_fd_sc_hd__o211a_1 _17476_ (.A1(_08870_),
    .A2(_10010_),
    .B1(_10011_),
    .C1(_09231_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_2 _17477_ (.A0(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[30] ),
    .A1(_10010_),
    .S(_08307_),
    .X(_10012_));
 sky130_fd_sc_hd__and2_4 _17478_ (.A(_09661_),
    .B(_10012_),
    .X(_10013_));
 sky130_fd_sc_hd__clkbuf_1 _17479_ (.A(_10013_),
    .X(_00587_));
 sky130_fd_sc_hd__and3_1 _17480_ (.A(_09990_),
    .B(_10000_),
    .C(_10008_),
    .X(_10014_));
 sky130_fd_sc_hd__nand2_1 _17481_ (.A(_09194_),
    .B(_09189_),
    .Y(_10015_));
 sky130_fd_sc_hd__a21o_1 _17482_ (.A1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[25] ),
    .A2(_10015_),
    .B1(_09418_),
    .X(_10016_));
 sky130_fd_sc_hd__a31o_1 _17483_ (.A1(_09625_),
    .A2(_09919_),
    .A3(_10016_),
    .B1(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[27] ),
    .X(_10017_));
 sky130_fd_sc_hd__xnor2_1 _17484_ (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[31] ),
    .B(_10005_),
    .Y(_10018_));
 sky130_fd_sc_hd__xnor2_1 _17485_ (.A(_10017_),
    .B(_10018_),
    .Y(_10019_));
 sky130_fd_sc_hd__o21ai_1 _17486_ (.A1(_10014_),
    .A2(_10019_),
    .B1(_05316_),
    .Y(_10020_));
 sky130_fd_sc_hd__a21o_1 _17487_ (.A1(_10014_),
    .A2(_10019_),
    .B1(_10020_),
    .X(_10021_));
 sky130_fd_sc_hd__o211a_1 _17488_ (.A1(net989),
    .A2(_08183_),
    .B1(_10021_),
    .C1(_09231_),
    .X(_00588_));
 sky130_fd_sc_hd__clkbuf_4 _17489_ (.A(\top_inst.grid_inst.data_path_wires[11][0] ),
    .X(_10022_));
 sky130_fd_sc_hd__or2_1 _17490_ (.A(_05736_),
    .B(_09187_),
    .X(_10023_));
 sky130_fd_sc_hd__buf_2 _17491_ (.A(_07617_),
    .X(_10024_));
 sky130_fd_sc_hd__o211a_1 _17492_ (.A1(_10022_),
    .A2(_07611_),
    .B1(_10023_),
    .C1(_10024_),
    .X(_00589_));
 sky130_fd_sc_hd__clkbuf_4 _17493_ (.A(\top_inst.grid_inst.data_path_wires[11][1] ),
    .X(_10025_));
 sky130_fd_sc_hd__or2_1 _17494_ (.A(_05736_),
    .B(_09192_),
    .X(_10026_));
 sky130_fd_sc_hd__o211a_1 _17495_ (.A1(_10025_),
    .A2(_07611_),
    .B1(_10026_),
    .C1(_10024_),
    .X(_00590_));
 sky130_fd_sc_hd__clkbuf_4 _17496_ (.A(\top_inst.grid_inst.data_path_wires[11][2] ),
    .X(_10027_));
 sky130_fd_sc_hd__or2_1 _17497_ (.A(_05736_),
    .B(_09197_),
    .X(_10028_));
 sky130_fd_sc_hd__o211a_1 _17498_ (.A1(_10027_),
    .A2(_07611_),
    .B1(_10028_),
    .C1(_10024_),
    .X(_00591_));
 sky130_fd_sc_hd__clkbuf_4 _17499_ (.A(\top_inst.grid_inst.data_path_wires[11][3] ),
    .X(_10029_));
 sky130_fd_sc_hd__buf_2 _17500_ (.A(_04858_),
    .X(_10030_));
 sky130_fd_sc_hd__or2_1 _17501_ (.A(_10030_),
    .B(_09202_),
    .X(_10031_));
 sky130_fd_sc_hd__o211a_1 _17502_ (.A1(_10029_),
    .A2(_07611_),
    .B1(_10031_),
    .C1(_10024_),
    .X(_00592_));
 sky130_fd_sc_hd__clkbuf_4 _17503_ (.A(\top_inst.grid_inst.data_path_wires[11][4] ),
    .X(_10032_));
 sky130_fd_sc_hd__clkbuf_4 _17504_ (.A(_04865_),
    .X(_10033_));
 sky130_fd_sc_hd__or2_1 _17505_ (.A(_10030_),
    .B(_09206_),
    .X(_10034_));
 sky130_fd_sc_hd__o211a_1 _17506_ (.A1(_10032_),
    .A2(_10033_),
    .B1(_10034_),
    .C1(_10024_),
    .X(_00593_));
 sky130_fd_sc_hd__clkbuf_4 _17507_ (.A(\top_inst.grid_inst.data_path_wires[11][5] ),
    .X(_10035_));
 sky130_fd_sc_hd__or2_1 _17508_ (.A(_10030_),
    .B(_09210_),
    .X(_10036_));
 sky130_fd_sc_hd__o211a_1 _17509_ (.A1(_10035_),
    .A2(_10033_),
    .B1(_10036_),
    .C1(_10024_),
    .X(_00594_));
 sky130_fd_sc_hd__buf_2 _17510_ (.A(\top_inst.grid_inst.data_path_wires[11][6] ),
    .X(_10037_));
 sky130_fd_sc_hd__clkbuf_4 _17511_ (.A(_10037_),
    .X(_10038_));
 sky130_fd_sc_hd__or2_2 _17512_ (.A(_10030_),
    .B(_09215_),
    .X(_10039_));
 sky130_fd_sc_hd__o211a_1 _17513_ (.A1(_10038_),
    .A2(_10033_),
    .B1(_10039_),
    .C1(_10024_),
    .X(_00595_));
 sky130_fd_sc_hd__buf_4 _17514_ (.A(\top_inst.grid_inst.data_path_wires[11][7] ),
    .X(_10040_));
 sky130_fd_sc_hd__or2_1 _17515_ (.A(_10030_),
    .B(_09219_),
    .X(_10041_));
 sky130_fd_sc_hd__o211a_1 _17516_ (.A1(_10040_),
    .A2(_10033_),
    .B1(_10041_),
    .C1(_10024_),
    .X(_00596_));
 sky130_fd_sc_hd__clkbuf_4 _17517_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[0] ),
    .X(_10042_));
 sky130_fd_sc_hd__or2_1 _17518_ (.A(_10042_),
    .B(_09199_),
    .X(_10043_));
 sky130_fd_sc_hd__o211a_1 _17519_ (.A1(_10022_),
    .A2(_08681_),
    .B1(_10043_),
    .C1(_10024_),
    .X(_00597_));
 sky130_fd_sc_hd__clkbuf_4 _17520_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[1] ),
    .X(_10044_));
 sky130_fd_sc_hd__or2_1 _17521_ (.A(_10044_),
    .B(_09199_),
    .X(_10045_));
 sky130_fd_sc_hd__o211a_1 _17522_ (.A1(_10025_),
    .A2(_08681_),
    .B1(_10045_),
    .C1(_10024_),
    .X(_00598_));
 sky130_fd_sc_hd__clkbuf_4 _17523_ (.A(_05755_),
    .X(_10046_));
 sky130_fd_sc_hd__clkbuf_4 _17524_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[2] ),
    .X(_10047_));
 sky130_fd_sc_hd__or2_1 _17525_ (.A(_10047_),
    .B(_09199_),
    .X(_10048_));
 sky130_fd_sc_hd__clkbuf_4 _17526_ (.A(_07617_),
    .X(_10049_));
 sky130_fd_sc_hd__o211a_1 _17527_ (.A1(_10027_),
    .A2(_10046_),
    .B1(_10048_),
    .C1(_10049_),
    .X(_00599_));
 sky130_fd_sc_hd__clkbuf_4 _17528_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[3] ),
    .X(_10050_));
 sky130_fd_sc_hd__or2_1 _17529_ (.A(_10050_),
    .B(_09199_),
    .X(_10051_));
 sky130_fd_sc_hd__o211a_1 _17530_ (.A1(_10029_),
    .A2(_10046_),
    .B1(_10051_),
    .C1(_10049_),
    .X(_00600_));
 sky130_fd_sc_hd__clkbuf_4 _17531_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[4] ),
    .X(_10052_));
 sky130_fd_sc_hd__or2_1 _17532_ (.A(_10052_),
    .B(_09199_),
    .X(_10053_));
 sky130_fd_sc_hd__o211a_1 _17533_ (.A1(_10032_),
    .A2(_10046_),
    .B1(_10053_),
    .C1(_10049_),
    .X(_00601_));
 sky130_fd_sc_hd__clkbuf_4 _17534_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[5] ),
    .X(_10054_));
 sky130_fd_sc_hd__or2_1 _17535_ (.A(_10054_),
    .B(_09199_),
    .X(_10055_));
 sky130_fd_sc_hd__o211a_1 _17536_ (.A1(_10035_),
    .A2(_10046_),
    .B1(_10055_),
    .C1(_10049_),
    .X(_00602_));
 sky130_fd_sc_hd__buf_2 _17537_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[6] ),
    .X(_10056_));
 sky130_fd_sc_hd__buf_2 _17538_ (.A(_05772_),
    .X(_10057_));
 sky130_fd_sc_hd__or2_1 _17539_ (.A(_10056_),
    .B(_10057_),
    .X(_10058_));
 sky130_fd_sc_hd__o211a_1 _17540_ (.A1(_10038_),
    .A2(_10046_),
    .B1(_10058_),
    .C1(_10049_),
    .X(_00603_));
 sky130_fd_sc_hd__clkbuf_4 _17541_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[7] ),
    .X(_10059_));
 sky130_fd_sc_hd__or2_1 _17542_ (.A(_10059_),
    .B(_10057_),
    .X(_10060_));
 sky130_fd_sc_hd__o211a_1 _17543_ (.A1(_10040_),
    .A2(_10046_),
    .B1(_10060_),
    .C1(_10049_),
    .X(_00604_));
 sky130_fd_sc_hd__and3_1 _17544_ (.A(_10022_),
    .B(_10042_),
    .C(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[0] ),
    .X(_10061_));
 sky130_fd_sc_hd__a21oi_1 _17545_ (.A1(_10022_),
    .A2(_10042_),
    .B1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[0] ),
    .Y(_10062_));
 sky130_fd_sc_hd__o21ai_1 _17546_ (.A1(_10061_),
    .A2(_10062_),
    .B1(_08181_),
    .Y(_10063_));
 sky130_fd_sc_hd__o211a_1 _17547_ (.A1(net1041),
    .A2(_08183_),
    .B1(_10063_),
    .C1(_10049_),
    .X(_00605_));
 sky130_fd_sc_hd__a22o_1 _17548_ (.A1(\top_inst.grid_inst.data_path_wires[11][0] ),
    .A2(_10044_),
    .B1(_10042_),
    .B2(_10025_),
    .X(_10064_));
 sky130_fd_sc_hd__nand4_2 _17549_ (.A(_10025_),
    .B(_10022_),
    .C(_10044_),
    .D(_10042_),
    .Y(_10065_));
 sky130_fd_sc_hd__nand3_1 _17550_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[1] ),
    .B(_10064_),
    .C(_10065_),
    .Y(_10066_));
 sky130_fd_sc_hd__a21o_1 _17551_ (.A1(_10064_),
    .A2(_10065_),
    .B1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[1] ),
    .X(_10067_));
 sky130_fd_sc_hd__a21o_1 _17552_ (.A1(_10066_),
    .A2(_10067_),
    .B1(_10061_),
    .X(_10068_));
 sky130_fd_sc_hd__nand3_2 _17553_ (.A(_10061_),
    .B(_10066_),
    .C(_10067_),
    .Y(_10069_));
 sky130_fd_sc_hd__a21o_1 _17554_ (.A1(_10068_),
    .A2(_10069_),
    .B1(_06682_),
    .X(_10070_));
 sky130_fd_sc_hd__o211a_1 _17555_ (.A1(net867),
    .A2(_08183_),
    .B1(_10070_),
    .C1(_10049_),
    .X(_00606_));
 sky130_fd_sc_hd__buf_4 _17556_ (.A(_05732_),
    .X(_10071_));
 sky130_fd_sc_hd__nand2_1 _17557_ (.A(_10022_),
    .B(_10047_),
    .Y(_10072_));
 sky130_fd_sc_hd__a22o_1 _17558_ (.A1(_10025_),
    .A2(_10044_),
    .B1(_10042_),
    .B2(_10027_),
    .X(_10073_));
 sky130_fd_sc_hd__nand4_1 _17559_ (.A(_10027_),
    .B(_10025_),
    .C(_10044_),
    .D(_10042_),
    .Y(_10074_));
 sky130_fd_sc_hd__nand2_1 _17560_ (.A(_10073_),
    .B(_10074_),
    .Y(_10075_));
 sky130_fd_sc_hd__xor2_1 _17561_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[2] ),
    .B(_10075_),
    .X(_10076_));
 sky130_fd_sc_hd__nand2_1 _17562_ (.A(_10065_),
    .B(_10066_),
    .Y(_10077_));
 sky130_fd_sc_hd__xor2_1 _17563_ (.A(_10076_),
    .B(_10077_),
    .X(_10078_));
 sky130_fd_sc_hd__or2_1 _17564_ (.A(_10072_),
    .B(_10078_),
    .X(_10079_));
 sky130_fd_sc_hd__nand2_1 _17565_ (.A(_10072_),
    .B(_10078_),
    .Y(_10080_));
 sky130_fd_sc_hd__and2_1 _17566_ (.A(_10079_),
    .B(_10080_),
    .X(_10081_));
 sky130_fd_sc_hd__xnor2_1 _17567_ (.A(_10069_),
    .B(_10081_),
    .Y(_10082_));
 sky130_fd_sc_hd__inv_2 _17568_ (.A(net1036),
    .Y(_10083_));
 sky130_fd_sc_hd__nand2_1 _17569_ (.A(_10083_),
    .B(_05403_),
    .Y(_10084_));
 sky130_fd_sc_hd__o211a_1 _17570_ (.A1(_10071_),
    .A2(_10082_),
    .B1(_10084_),
    .C1(_10049_),
    .X(_00607_));
 sky130_fd_sc_hd__or2b_1 _17571_ (.A(_10069_),
    .B_N(_10081_),
    .X(_10085_));
 sky130_fd_sc_hd__or2b_1 _17572_ (.A(_10076_),
    .B_N(_10077_),
    .X(_10086_));
 sky130_fd_sc_hd__a22o_1 _17573_ (.A1(_10022_),
    .A2(_10050_),
    .B1(_10047_),
    .B2(_10025_),
    .X(_10087_));
 sky130_fd_sc_hd__and3_1 _17574_ (.A(\top_inst.grid_inst.data_path_wires[11][1] ),
    .B(\top_inst.grid_inst.data_path_wires[11][0] ),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[3] ),
    .X(_10088_));
 sky130_fd_sc_hd__nand2_2 _17575_ (.A(_10047_),
    .B(_10088_),
    .Y(_10089_));
 sky130_fd_sc_hd__nand2_1 _17576_ (.A(_10087_),
    .B(_10089_),
    .Y(_10090_));
 sky130_fd_sc_hd__a22o_1 _17577_ (.A1(_10027_),
    .A2(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[0] ),
    .B2(_10029_),
    .X(_10091_));
 sky130_fd_sc_hd__nand4_1 _17578_ (.A(_10029_),
    .B(_10027_),
    .C(_10044_),
    .D(_10042_),
    .Y(_10092_));
 sky130_fd_sc_hd__and3_1 _17579_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[3] ),
    .B(_10091_),
    .C(_10092_),
    .X(_10093_));
 sky130_fd_sc_hd__a21oi_1 _17580_ (.A1(_10091_),
    .A2(_10092_),
    .B1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[3] ),
    .Y(_10094_));
 sky130_fd_sc_hd__or2_1 _17581_ (.A(_10093_),
    .B(_10094_),
    .X(_10095_));
 sky130_fd_sc_hd__a21boi_2 _17582_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[2] ),
    .A2(_10073_),
    .B1_N(_10074_),
    .Y(_10096_));
 sky130_fd_sc_hd__xnor2_1 _17583_ (.A(_10095_),
    .B(_10096_),
    .Y(_10097_));
 sky130_fd_sc_hd__xnor2_1 _17584_ (.A(_10090_),
    .B(_10097_),
    .Y(_10098_));
 sky130_fd_sc_hd__a21o_1 _17585_ (.A1(_10086_),
    .A2(_10079_),
    .B1(_10098_),
    .X(_10099_));
 sky130_fd_sc_hd__inv_2 _17586_ (.A(_10099_),
    .Y(_10100_));
 sky130_fd_sc_hd__and3_1 _17587_ (.A(_10086_),
    .B(_10079_),
    .C(_10098_),
    .X(_10101_));
 sky130_fd_sc_hd__or3_1 _17588_ (.A(_10085_),
    .B(_10100_),
    .C(_10101_),
    .X(_10102_));
 sky130_fd_sc_hd__o21ai_1 _17589_ (.A1(_10100_),
    .A2(_10101_),
    .B1(_10085_),
    .Y(_10103_));
 sky130_fd_sc_hd__and2_1 _17590_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[3] ),
    .B(_05730_),
    .X(_10104_));
 sky130_fd_sc_hd__a31o_1 _17591_ (.A1(_05887_),
    .A2(_10102_),
    .A3(_10103_),
    .B1(_10104_),
    .X(_10105_));
 sky130_fd_sc_hd__and2_1 _17592_ (.A(_09661_),
    .B(_10105_),
    .X(_10106_));
 sky130_fd_sc_hd__clkbuf_1 _17593_ (.A(_10106_),
    .X(_00608_));
 sky130_fd_sc_hd__a22o_1 _17594_ (.A1(\top_inst.grid_inst.data_path_wires[11][3] ),
    .A2(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[11][4] ),
    .X(_10107_));
 sky130_fd_sc_hd__nand4_1 _17595_ (.A(_10032_),
    .B(_10029_),
    .C(_10044_),
    .D(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[0] ),
    .Y(_10108_));
 sky130_fd_sc_hd__nand2_1 _17596_ (.A(_10107_),
    .B(_10108_),
    .Y(_10109_));
 sky130_fd_sc_hd__xor2_2 _17597_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[4] ),
    .B(_10109_),
    .X(_10110_));
 sky130_fd_sc_hd__xor2_2 _17598_ (.A(_10089_),
    .B(_10110_),
    .X(_10111_));
 sky130_fd_sc_hd__a21bo_1 _17599_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[3] ),
    .A2(_10091_),
    .B1_N(_10092_),
    .X(_10112_));
 sky130_fd_sc_hd__xnor2_2 _17600_ (.A(_10111_),
    .B(_10112_),
    .Y(_10113_));
 sky130_fd_sc_hd__nand2_1 _17601_ (.A(_10027_),
    .B(_10047_),
    .Y(_10114_));
 sky130_fd_sc_hd__a22o_1 _17602_ (.A1(\top_inst.grid_inst.data_path_wires[11][0] ),
    .A2(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[11][1] ),
    .X(_10115_));
 sky130_fd_sc_hd__a21bo_1 _17603_ (.A1(_10052_),
    .A2(_10088_),
    .B1_N(_10115_),
    .X(_10116_));
 sky130_fd_sc_hd__xor2_2 _17604_ (.A(_10114_),
    .B(_10116_),
    .X(_10117_));
 sky130_fd_sc_hd__xor2_2 _17605_ (.A(_10113_),
    .B(_10117_),
    .X(_10118_));
 sky130_fd_sc_hd__or2_1 _17606_ (.A(_10090_),
    .B(_10097_),
    .X(_10119_));
 sky130_fd_sc_hd__o21ai_2 _17607_ (.A1(_10095_),
    .A2(_10096_),
    .B1(_10119_),
    .Y(_10120_));
 sky130_fd_sc_hd__xor2_2 _17608_ (.A(_10118_),
    .B(_10120_),
    .X(_10121_));
 sky130_fd_sc_hd__nand2_1 _17609_ (.A(_10099_),
    .B(_10102_),
    .Y(_10122_));
 sky130_fd_sc_hd__nor2_1 _17610_ (.A(_10121_),
    .B(_10122_),
    .Y(_10123_));
 sky130_fd_sc_hd__a21o_1 _17611_ (.A1(_10121_),
    .A2(_10122_),
    .B1(_09292_),
    .X(_10124_));
 sky130_fd_sc_hd__o221a_1 _17612_ (.A1(net1053),
    .A2(_09266_),
    .B1(_10123_),
    .B2(_10124_),
    .C1(_09886_),
    .X(_00609_));
 sky130_fd_sc_hd__nor2_1 _17613_ (.A(_10102_),
    .B(_10121_),
    .Y(_10125_));
 sky130_fd_sc_hd__and2b_1 _17614_ (.A_N(_10113_),
    .B(_10117_),
    .X(_10126_));
 sky130_fd_sc_hd__nand2_1 _17615_ (.A(_10022_),
    .B(_10054_),
    .Y(_10127_));
 sky130_fd_sc_hd__nand2_1 _17616_ (.A(_10029_),
    .B(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[2] ),
    .Y(_10128_));
 sky130_fd_sc_hd__and3_1 _17617_ (.A(\top_inst.grid_inst.data_path_wires[11][2] ),
    .B(\top_inst.grid_inst.data_path_wires[11][1] ),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[4] ),
    .X(_10129_));
 sky130_fd_sc_hd__a22o_1 _17618_ (.A1(\top_inst.grid_inst.data_path_wires[11][1] ),
    .A2(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[11][2] ),
    .X(_10130_));
 sky130_fd_sc_hd__a21bo_1 _17619_ (.A1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[3] ),
    .A2(_10129_),
    .B1_N(_10130_),
    .X(_10131_));
 sky130_fd_sc_hd__xor2_2 _17620_ (.A(_10128_),
    .B(_10131_),
    .X(_10132_));
 sky130_fd_sc_hd__xnor2_2 _17621_ (.A(_10127_),
    .B(_10132_),
    .Y(_10133_));
 sky130_fd_sc_hd__a21boi_2 _17622_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[4] ),
    .A2(_10107_),
    .B1_N(_10108_),
    .Y(_10134_));
 sky130_fd_sc_hd__a32o_1 _17623_ (.A1(_10027_),
    .A2(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[2] ),
    .A3(_10115_),
    .B1(_10088_),
    .B2(_10052_),
    .X(_10135_));
 sky130_fd_sc_hd__a22o_1 _17624_ (.A1(\top_inst.grid_inst.data_path_wires[11][4] ),
    .A2(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[11][5] ),
    .X(_10136_));
 sky130_fd_sc_hd__nand4_1 _17625_ (.A(\top_inst.grid_inst.data_path_wires[11][5] ),
    .B(\top_inst.grid_inst.data_path_wires[11][4] ),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[0] ),
    .Y(_10137_));
 sky130_fd_sc_hd__nand2_1 _17626_ (.A(_10136_),
    .B(_10137_),
    .Y(_10138_));
 sky130_fd_sc_hd__xor2_2 _17627_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[5] ),
    .B(_10138_),
    .X(_10139_));
 sky130_fd_sc_hd__xnor2_1 _17628_ (.A(_10135_),
    .B(_10139_),
    .Y(_10140_));
 sky130_fd_sc_hd__xnor2_2 _17629_ (.A(_10134_),
    .B(_10140_),
    .Y(_10141_));
 sky130_fd_sc_hd__xor2_2 _17630_ (.A(_10133_),
    .B(_10141_),
    .X(_10142_));
 sky130_fd_sc_hd__xor2_2 _17631_ (.A(_10126_),
    .B(_10142_),
    .X(_10143_));
 sky130_fd_sc_hd__nor2_1 _17632_ (.A(_10089_),
    .B(_10110_),
    .Y(_10144_));
 sky130_fd_sc_hd__a21o_1 _17633_ (.A1(_10111_),
    .A2(_10112_),
    .B1(_10144_),
    .X(_10145_));
 sky130_fd_sc_hd__xnor2_2 _17634_ (.A(_10143_),
    .B(_10145_),
    .Y(_10146_));
 sky130_fd_sc_hd__or2b_1 _17635_ (.A(_10118_),
    .B_N(_10120_),
    .X(_10147_));
 sky130_fd_sc_hd__o21a_1 _17636_ (.A1(_10099_),
    .A2(_10121_),
    .B1(_10147_),
    .X(_10148_));
 sky130_fd_sc_hd__xor2_1 _17637_ (.A(_10146_),
    .B(_10148_),
    .X(_10149_));
 sky130_fd_sc_hd__nand2_1 _17638_ (.A(_10125_),
    .B(_10149_),
    .Y(_10150_));
 sky130_fd_sc_hd__o21a_1 _17639_ (.A1(_10125_),
    .A2(_10149_),
    .B1(_08265_),
    .X(_10151_));
 sky130_fd_sc_hd__a22o_1 _17640_ (.A1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[5] ),
    .A2(_09496_),
    .B1(_10150_),
    .B2(_10151_),
    .X(_10152_));
 sky130_fd_sc_hd__and2_1 _17641_ (.A(_09661_),
    .B(_10152_),
    .X(_10153_));
 sky130_fd_sc_hd__clkbuf_1 _17642_ (.A(_10153_),
    .X(_00610_));
 sky130_fd_sc_hd__nand2_1 _17643_ (.A(_10126_),
    .B(_10142_),
    .Y(_10154_));
 sky130_fd_sc_hd__nand2_1 _17644_ (.A(_10143_),
    .B(_10145_),
    .Y(_10155_));
 sky130_fd_sc_hd__or2b_1 _17645_ (.A(_10139_),
    .B_N(_10135_),
    .X(_10156_));
 sky130_fd_sc_hd__or2b_1 _17646_ (.A(_10134_),
    .B_N(_10140_),
    .X(_10157_));
 sky130_fd_sc_hd__and2_1 _17647_ (.A(_10133_),
    .B(_10141_),
    .X(_10158_));
 sky130_fd_sc_hd__a21boi_1 _17648_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[5] ),
    .A2(_10136_),
    .B1_N(_10137_),
    .Y(_10159_));
 sky130_fd_sc_hd__o2bb2a_1 _17649_ (.A1_N(_10050_),
    .A2_N(_10129_),
    .B1(_10131_),
    .B2(_10128_),
    .X(_10160_));
 sky130_fd_sc_hd__a22o_1 _17650_ (.A1(\top_inst.grid_inst.data_path_wires[11][5] ),
    .A2(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[0] ),
    .B2(_10037_),
    .X(_10161_));
 sky130_fd_sc_hd__nand4_1 _17651_ (.A(_10037_),
    .B(\top_inst.grid_inst.data_path_wires[11][5] ),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[0] ),
    .Y(_10162_));
 sky130_fd_sc_hd__nand2_1 _17652_ (.A(_10161_),
    .B(_10162_),
    .Y(_10163_));
 sky130_fd_sc_hd__xor2_2 _17653_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[6] ),
    .B(_10163_),
    .X(_10164_));
 sky130_fd_sc_hd__xor2_1 _17654_ (.A(_10160_),
    .B(_10164_),
    .X(_10165_));
 sky130_fd_sc_hd__xnor2_1 _17655_ (.A(_10159_),
    .B(_10165_),
    .Y(_10166_));
 sky130_fd_sc_hd__or2b_1 _17656_ (.A(_10127_),
    .B_N(_10132_),
    .X(_10167_));
 sky130_fd_sc_hd__a22oi_1 _17657_ (.A1(_10022_),
    .A2(_10056_),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[5] ),
    .B2(_10025_),
    .Y(_10168_));
 sky130_fd_sc_hd__and4_1 _17658_ (.A(\top_inst.grid_inst.data_path_wires[11][1] ),
    .B(\top_inst.grid_inst.data_path_wires[11][0] ),
    .C(_10056_),
    .D(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[5] ),
    .X(_10169_));
 sky130_fd_sc_hd__nor2_1 _17659_ (.A(_10168_),
    .B(_10169_),
    .Y(_10170_));
 sky130_fd_sc_hd__a22oi_1 _17660_ (.A1(\top_inst.grid_inst.data_path_wires[11][2] ),
    .A2(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[11][3] ),
    .Y(_10171_));
 sky130_fd_sc_hd__and4_1 _17661_ (.A(\top_inst.grid_inst.data_path_wires[11][3] ),
    .B(\top_inst.grid_inst.data_path_wires[11][2] ),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[3] ),
    .X(_10172_));
 sky130_fd_sc_hd__and4bb_1 _17662_ (.A_N(_10171_),
    .B_N(_10172_),
    .C(_10032_),
    .D(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[2] ),
    .X(_10173_));
 sky130_fd_sc_hd__o2bb2a_1 _17663_ (.A1_N(_10032_),
    .A2_N(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[2] ),
    .B1(_10171_),
    .B2(_10172_),
    .X(_10174_));
 sky130_fd_sc_hd__nor2_1 _17664_ (.A(_10173_),
    .B(_10174_),
    .Y(_10175_));
 sky130_fd_sc_hd__xnor2_1 _17665_ (.A(_10170_),
    .B(_10175_),
    .Y(_10176_));
 sky130_fd_sc_hd__xor2_1 _17666_ (.A(_10167_),
    .B(_10176_),
    .X(_10177_));
 sky130_fd_sc_hd__nand2_1 _17667_ (.A(_10166_),
    .B(_10177_),
    .Y(_10178_));
 sky130_fd_sc_hd__or2_1 _17668_ (.A(_10166_),
    .B(_10177_),
    .X(_10179_));
 sky130_fd_sc_hd__and3_1 _17669_ (.A(_10158_),
    .B(_10178_),
    .C(_10179_),
    .X(_10180_));
 sky130_fd_sc_hd__a21oi_1 _17670_ (.A1(_10178_),
    .A2(_10179_),
    .B1(_10158_),
    .Y(_10181_));
 sky130_fd_sc_hd__a211oi_2 _17671_ (.A1(_10156_),
    .A2(_10157_),
    .B1(_10180_),
    .C1(_10181_),
    .Y(_10182_));
 sky130_fd_sc_hd__o211a_1 _17672_ (.A1(_10180_),
    .A2(_10181_),
    .B1(_10156_),
    .C1(_10157_),
    .X(_10183_));
 sky130_fd_sc_hd__a211o_1 _17673_ (.A1(_10154_),
    .A2(_10155_),
    .B1(_10182_),
    .C1(_10183_),
    .X(_10184_));
 sky130_fd_sc_hd__o211ai_1 _17674_ (.A1(_10182_),
    .A2(_10183_),
    .B1(_10154_),
    .C1(_10155_),
    .Y(_10185_));
 sky130_fd_sc_hd__and4bb_1 _17675_ (.A_N(_10147_),
    .B_N(_10146_),
    .C(_10184_),
    .D(_10185_),
    .X(_10186_));
 sky130_fd_sc_hd__o2bb2a_1 _17676_ (.A1_N(_10184_),
    .A2_N(_10185_),
    .B1(_10147_),
    .B2(_10146_),
    .X(_10187_));
 sky130_fd_sc_hd__nor2_1 _17677_ (.A(_10186_),
    .B(_10187_),
    .Y(_10188_));
 sky130_fd_sc_hd__o31a_1 _17678_ (.A1(_10099_),
    .A2(_10121_),
    .A3(_10146_),
    .B1(_10150_),
    .X(_10189_));
 sky130_fd_sc_hd__xnor2_1 _17679_ (.A(_10188_),
    .B(_10189_),
    .Y(_10190_));
 sky130_fd_sc_hd__mux2_1 _17680_ (.A0(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[6] ),
    .A1(_10190_),
    .S(_08307_),
    .X(_10191_));
 sky130_fd_sc_hd__and2_1 _17681_ (.A(_09661_),
    .B(_10191_),
    .X(_10192_));
 sky130_fd_sc_hd__clkbuf_1 _17682_ (.A(_10192_),
    .X(_00611_));
 sky130_fd_sc_hd__or2b_1 _17683_ (.A(_10159_),
    .B_N(_10165_),
    .X(_10193_));
 sky130_fd_sc_hd__o21ai_2 _17684_ (.A1(_10160_),
    .A2(_10164_),
    .B1(_10193_),
    .Y(_10194_));
 sky130_fd_sc_hd__o21ai_1 _17685_ (.A1(_10167_),
    .A2(_10176_),
    .B1(_10178_),
    .Y(_10195_));
 sky130_fd_sc_hd__a21bo_1 _17686_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[6] ),
    .A2(_10161_),
    .B1_N(_10162_),
    .X(_10196_));
 sky130_fd_sc_hd__nor2_1 _17687_ (.A(_10172_),
    .B(_10173_),
    .Y(_10197_));
 sky130_fd_sc_hd__a22o_1 _17688_ (.A1(_10037_),
    .A2(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[11][7] ),
    .X(_10198_));
 sky130_fd_sc_hd__nand4_1 _17689_ (.A(\top_inst.grid_inst.data_path_wires[11][7] ),
    .B(_10037_),
    .C(_10044_),
    .D(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[0] ),
    .Y(_10199_));
 sky130_fd_sc_hd__nand2_1 _17690_ (.A(_10198_),
    .B(_10199_),
    .Y(_10200_));
 sky130_fd_sc_hd__xor2_2 _17691_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[7] ),
    .B(_10200_),
    .X(_10201_));
 sky130_fd_sc_hd__xor2_2 _17692_ (.A(_10197_),
    .B(_10201_),
    .X(_10202_));
 sky130_fd_sc_hd__xnor2_2 _17693_ (.A(_10196_),
    .B(_10202_),
    .Y(_10203_));
 sky130_fd_sc_hd__and2_1 _17694_ (.A(_10170_),
    .B(_10175_),
    .X(_10204_));
 sky130_fd_sc_hd__a22o_1 _17695_ (.A1(\top_inst.grid_inst.data_path_wires[11][3] ),
    .A2(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[11][4] ),
    .X(_10205_));
 sky130_fd_sc_hd__nand4_2 _17696_ (.A(_10032_),
    .B(_10029_),
    .C(_10052_),
    .D(_10050_),
    .Y(_10206_));
 sky130_fd_sc_hd__a22o_1 _17697_ (.A1(_10035_),
    .A2(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[2] ),
    .B1(_10205_),
    .B2(_10206_),
    .X(_10207_));
 sky130_fd_sc_hd__nand4_1 _17698_ (.A(_10035_),
    .B(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[2] ),
    .C(_10205_),
    .D(_10206_),
    .Y(_10208_));
 sky130_fd_sc_hd__nand2_1 _17699_ (.A(_10207_),
    .B(_10208_),
    .Y(_10209_));
 sky130_fd_sc_hd__nand2_1 _17700_ (.A(\top_inst.grid_inst.data_path_wires[11][2] ),
    .B(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[5] ),
    .Y(_10210_));
 sky130_fd_sc_hd__nand2_1 _17701_ (.A(\top_inst.grid_inst.data_path_wires[11][1] ),
    .B(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[6] ),
    .Y(_10211_));
 sky130_fd_sc_hd__and2b_1 _17702_ (.A_N(\top_inst.grid_inst.data_path_wires[11][0] ),
    .B(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[7] ),
    .X(_10212_));
 sky130_fd_sc_hd__xnor2_1 _17703_ (.A(_10211_),
    .B(_10212_),
    .Y(_10213_));
 sky130_fd_sc_hd__xnor2_1 _17704_ (.A(_10210_),
    .B(_10213_),
    .Y(_10214_));
 sky130_fd_sc_hd__xnor2_1 _17705_ (.A(_10169_),
    .B(_10214_),
    .Y(_10215_));
 sky130_fd_sc_hd__xor2_1 _17706_ (.A(_10209_),
    .B(_10215_),
    .X(_10216_));
 sky130_fd_sc_hd__xnor2_1 _17707_ (.A(_10204_),
    .B(_10216_),
    .Y(_10217_));
 sky130_fd_sc_hd__xnor2_1 _17708_ (.A(_10203_),
    .B(_10217_),
    .Y(_10218_));
 sky130_fd_sc_hd__xor2_1 _17709_ (.A(_10195_),
    .B(_10218_),
    .X(_10219_));
 sky130_fd_sc_hd__xnor2_1 _17710_ (.A(_10194_),
    .B(_10219_),
    .Y(_10220_));
 sky130_fd_sc_hd__nor2_1 _17711_ (.A(_10180_),
    .B(_10182_),
    .Y(_10221_));
 sky130_fd_sc_hd__xnor2_1 _17712_ (.A(_10220_),
    .B(_10221_),
    .Y(_10222_));
 sky130_fd_sc_hd__xnor2_1 _17713_ (.A(_10059_),
    .B(_10222_),
    .Y(_10223_));
 sky130_fd_sc_hd__xor2_1 _17714_ (.A(_10184_),
    .B(_10223_),
    .X(_10224_));
 sky130_fd_sc_hd__o21bai_2 _17715_ (.A1(_10187_),
    .A2(_10189_),
    .B1_N(_10186_),
    .Y(_10225_));
 sky130_fd_sc_hd__nor2_1 _17716_ (.A(_10224_),
    .B(_10225_),
    .Y(_10226_));
 sky130_fd_sc_hd__a21o_1 _17717_ (.A1(_10224_),
    .A2(_10225_),
    .B1(_05353_),
    .X(_10227_));
 sky130_fd_sc_hd__a2bb2o_1 _17718_ (.A1_N(_10226_),
    .A2_N(_10227_),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[7] ),
    .B2(_07816_),
    .X(_10228_));
 sky130_fd_sc_hd__and2_1 _17719_ (.A(_09661_),
    .B(_10228_),
    .X(_10229_));
 sky130_fd_sc_hd__clkbuf_1 _17720_ (.A(_10229_),
    .X(_00612_));
 sky130_fd_sc_hd__nor2_1 _17721_ (.A(_10197_),
    .B(_10201_),
    .Y(_10230_));
 sky130_fd_sc_hd__a21o_1 _17722_ (.A1(_10196_),
    .A2(_10202_),
    .B1(_10230_),
    .X(_10231_));
 sky130_fd_sc_hd__a21boi_2 _17723_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[7] ),
    .A2(_10198_),
    .B1_N(_10199_),
    .Y(_10232_));
 sky130_fd_sc_hd__nand2_1 _17724_ (.A(_10206_),
    .B(_10208_),
    .Y(_10233_));
 sky130_fd_sc_hd__o21ai_2 _17725_ (.A1(_10044_),
    .A2(_10042_),
    .B1(\top_inst.grid_inst.data_path_wires[11][7] ),
    .Y(_10234_));
 sky130_fd_sc_hd__and3_1 _17726_ (.A(\top_inst.grid_inst.data_path_wires[11][7] ),
    .B(_10044_),
    .C(_10042_),
    .X(_10235_));
 sky130_fd_sc_hd__nor2_4 _17727_ (.A(_10234_),
    .B(_10235_),
    .Y(_10236_));
 sky130_fd_sc_hd__xnor2_2 _17728_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[8] ),
    .B(_10236_),
    .Y(_10237_));
 sky130_fd_sc_hd__xnor2_2 _17729_ (.A(_10233_),
    .B(_10237_),
    .Y(_10238_));
 sky130_fd_sc_hd__xnor2_2 _17730_ (.A(_10232_),
    .B(_10238_),
    .Y(_10239_));
 sky130_fd_sc_hd__a22o_1 _17731_ (.A1(_10032_),
    .A2(_10052_),
    .B1(_10050_),
    .B2(_10035_),
    .X(_10240_));
 sky130_fd_sc_hd__nand4_2 _17732_ (.A(_10035_),
    .B(_10032_),
    .C(_10052_),
    .D(_10050_),
    .Y(_10241_));
 sky130_fd_sc_hd__a22o_1 _17733_ (.A1(_10038_),
    .A2(_10047_),
    .B1(_10240_),
    .B2(_10241_),
    .X(_10242_));
 sky130_fd_sc_hd__nand4_1 _17734_ (.A(_10038_),
    .B(_10047_),
    .C(_10240_),
    .D(_10241_),
    .Y(_10243_));
 sky130_fd_sc_hd__nand2_1 _17735_ (.A(_10242_),
    .B(_10243_),
    .Y(_10244_));
 sky130_fd_sc_hd__nand2_1 _17736_ (.A(_10029_),
    .B(_10054_),
    .Y(_10245_));
 sky130_fd_sc_hd__inv_2 _17737_ (.A(\top_inst.grid_inst.data_path_wires[11][1] ),
    .Y(_10246_));
 sky130_fd_sc_hd__and4_1 _17738_ (.A(\top_inst.grid_inst.data_path_wires[11][2] ),
    .B(_10246_),
    .C(_10059_),
    .D(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[6] ),
    .X(_10247_));
 sky130_fd_sc_hd__a22o_1 _17739_ (.A1(_10246_),
    .A2(_10059_),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[6] ),
    .B2(\top_inst.grid_inst.data_path_wires[11][2] ),
    .X(_10248_));
 sky130_fd_sc_hd__and2b_1 _17740_ (.A_N(_10247_),
    .B(_10248_),
    .X(_10249_));
 sky130_fd_sc_hd__xnor2_1 _17741_ (.A(_10245_),
    .B(_10249_),
    .Y(_10250_));
 sky130_fd_sc_hd__and3_1 _17742_ (.A(_10025_),
    .B(_10056_),
    .C(_10212_),
    .X(_10251_));
 sky130_fd_sc_hd__a31oi_2 _17743_ (.A1(_10027_),
    .A2(_10054_),
    .A3(_10213_),
    .B1(_10251_),
    .Y(_10252_));
 sky130_fd_sc_hd__xnor2_1 _17744_ (.A(_10250_),
    .B(_10252_),
    .Y(_10253_));
 sky130_fd_sc_hd__xnor2_1 _17745_ (.A(_10244_),
    .B(_10253_),
    .Y(_10254_));
 sky130_fd_sc_hd__nand2_1 _17746_ (.A(_10169_),
    .B(_10214_),
    .Y(_10255_));
 sky130_fd_sc_hd__o21a_1 _17747_ (.A1(_10209_),
    .A2(_10215_),
    .B1(_10255_),
    .X(_10256_));
 sky130_fd_sc_hd__xnor2_1 _17748_ (.A(_10254_),
    .B(_10256_),
    .Y(_10257_));
 sky130_fd_sc_hd__xnor2_1 _17749_ (.A(_10239_),
    .B(_10257_),
    .Y(_10258_));
 sky130_fd_sc_hd__nand2_1 _17750_ (.A(_10204_),
    .B(_10216_),
    .Y(_10259_));
 sky130_fd_sc_hd__o21a_1 _17751_ (.A1(_10203_),
    .A2(_10217_),
    .B1(_10259_),
    .X(_10260_));
 sky130_fd_sc_hd__xor2_1 _17752_ (.A(_10258_),
    .B(_10260_),
    .X(_10261_));
 sky130_fd_sc_hd__xnor2_1 _17753_ (.A(_10231_),
    .B(_10261_),
    .Y(_10262_));
 sky130_fd_sc_hd__or2b_1 _17754_ (.A(_10218_),
    .B_N(_10195_),
    .X(_10263_));
 sky130_fd_sc_hd__or2b_1 _17755_ (.A(_10219_),
    .B_N(_10194_),
    .X(_10264_));
 sky130_fd_sc_hd__and2_1 _17756_ (.A(_10263_),
    .B(_10264_),
    .X(_10265_));
 sky130_fd_sc_hd__xnor2_1 _17757_ (.A(_10262_),
    .B(_10265_),
    .Y(_10266_));
 sky130_fd_sc_hd__and2b_1 _17758_ (.A_N(_10221_),
    .B(_10220_),
    .X(_10267_));
 sky130_fd_sc_hd__a21oi_1 _17759_ (.A1(_10059_),
    .A2(_10222_),
    .B1(_10267_),
    .Y(_10268_));
 sky130_fd_sc_hd__nor2_1 _17760_ (.A(_10266_),
    .B(_10268_),
    .Y(_10269_));
 sky130_fd_sc_hd__and2_1 _17761_ (.A(_10266_),
    .B(_10268_),
    .X(_10270_));
 sky130_fd_sc_hd__nor2_1 _17762_ (.A(_10269_),
    .B(_10270_),
    .Y(_10271_));
 sky130_fd_sc_hd__nor2_1 _17763_ (.A(_10184_),
    .B(_10223_),
    .Y(_10272_));
 sky130_fd_sc_hd__a21o_1 _17764_ (.A1(_10224_),
    .A2(_10225_),
    .B1(_10272_),
    .X(_10273_));
 sky130_fd_sc_hd__nand2_1 _17765_ (.A(_10271_),
    .B(_10273_),
    .Y(_10274_));
 sky130_fd_sc_hd__o21a_1 _17766_ (.A1(_10271_),
    .A2(_10273_),
    .B1(_08265_),
    .X(_10275_));
 sky130_fd_sc_hd__a22o_1 _17767_ (.A1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[8] ),
    .A2(_09496_),
    .B1(_10274_),
    .B2(_10275_),
    .X(_10276_));
 sky130_fd_sc_hd__and2_1 _17768_ (.A(_09661_),
    .B(_10276_),
    .X(_10277_));
 sky130_fd_sc_hd__clkbuf_1 _17769_ (.A(_10277_),
    .X(_00613_));
 sky130_fd_sc_hd__nor2_1 _17770_ (.A(_10262_),
    .B(_10265_),
    .Y(_10278_));
 sky130_fd_sc_hd__a21o_1 _17771_ (.A1(_10271_),
    .A2(_10273_),
    .B1(_10269_),
    .X(_10279_));
 sky130_fd_sc_hd__or2b_1 _17772_ (.A(_10237_),
    .B_N(_10233_),
    .X(_10280_));
 sky130_fd_sc_hd__or2b_1 _17773_ (.A(_10232_),
    .B_N(_10238_),
    .X(_10281_));
 sky130_fd_sc_hd__nand2_1 _17774_ (.A(_10280_),
    .B(_10281_),
    .Y(_10282_));
 sky130_fd_sc_hd__clkbuf_4 _17775_ (.A(_10235_),
    .X(_10283_));
 sky130_fd_sc_hd__a21o_1 _17776_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[8] ),
    .A2(_10236_),
    .B1(_10283_),
    .X(_10284_));
 sky130_fd_sc_hd__xnor2_1 _17777_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[9] ),
    .B(_10236_),
    .Y(_10285_));
 sky130_fd_sc_hd__a21oi_1 _17778_ (.A1(_10241_),
    .A2(_10243_),
    .B1(_10285_),
    .Y(_10286_));
 sky130_fd_sc_hd__and3_1 _17779_ (.A(_10241_),
    .B(_10243_),
    .C(_10285_),
    .X(_10287_));
 sky130_fd_sc_hd__nor2_1 _17780_ (.A(_10286_),
    .B(_10287_),
    .Y(_10288_));
 sky130_fd_sc_hd__xor2_1 _17781_ (.A(_10284_),
    .B(_10288_),
    .X(_10289_));
 sky130_fd_sc_hd__or2b_1 _17782_ (.A(_10252_),
    .B_N(_10250_),
    .X(_10290_));
 sky130_fd_sc_hd__or2b_1 _17783_ (.A(_10244_),
    .B_N(_10253_),
    .X(_10291_));
 sky130_fd_sc_hd__a22o_1 _17784_ (.A1(\top_inst.grid_inst.data_path_wires[11][5] ),
    .A2(_10052_),
    .B1(_10050_),
    .B2(_10037_),
    .X(_10292_));
 sky130_fd_sc_hd__and4_1 _17785_ (.A(\top_inst.grid_inst.data_path_wires[11][6] ),
    .B(\top_inst.grid_inst.data_path_wires[11][5] ),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[3] ),
    .X(_10293_));
 sky130_fd_sc_hd__inv_2 _17786_ (.A(_10293_),
    .Y(_10294_));
 sky130_fd_sc_hd__and2_1 _17787_ (.A(_10292_),
    .B(_10294_),
    .X(_10295_));
 sky130_fd_sc_hd__nand2_4 _17788_ (.A(_10040_),
    .B(_10047_),
    .Y(_10296_));
 sky130_fd_sc_hd__xor2_1 _17789_ (.A(_10295_),
    .B(_10296_),
    .X(_10297_));
 sky130_fd_sc_hd__nand2_1 _17790_ (.A(_10032_),
    .B(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[5] ),
    .Y(_10298_));
 sky130_fd_sc_hd__and4b_1 _17791_ (.A_N(\top_inst.grid_inst.data_path_wires[11][2] ),
    .B(_10059_),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[6] ),
    .D(\top_inst.grid_inst.data_path_wires[11][3] ),
    .X(_10299_));
 sky130_fd_sc_hd__inv_2 _17792_ (.A(_10059_),
    .Y(_10300_));
 sky130_fd_sc_hd__o2bb2a_1 _17793_ (.A1_N(\top_inst.grid_inst.data_path_wires[11][3] ),
    .A2_N(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[6] ),
    .B1(_10300_),
    .B2(\top_inst.grid_inst.data_path_wires[11][2] ),
    .X(_10301_));
 sky130_fd_sc_hd__nor2_1 _17794_ (.A(_10299_),
    .B(_10301_),
    .Y(_10302_));
 sky130_fd_sc_hd__xnor2_1 _17795_ (.A(_10298_),
    .B(_10302_),
    .Y(_10303_));
 sky130_fd_sc_hd__a31oi_2 _17796_ (.A1(_10029_),
    .A2(_10054_),
    .A3(_10248_),
    .B1(_10247_),
    .Y(_10304_));
 sky130_fd_sc_hd__xnor2_1 _17797_ (.A(_10303_),
    .B(_10304_),
    .Y(_10305_));
 sky130_fd_sc_hd__xor2_1 _17798_ (.A(_10297_),
    .B(_10305_),
    .X(_10306_));
 sky130_fd_sc_hd__a21oi_1 _17799_ (.A1(_10290_),
    .A2(_10291_),
    .B1(_10306_),
    .Y(_10307_));
 sky130_fd_sc_hd__and3_1 _17800_ (.A(_10290_),
    .B(_10291_),
    .C(_10306_),
    .X(_10308_));
 sky130_fd_sc_hd__nor2_1 _17801_ (.A(_10307_),
    .B(_10308_),
    .Y(_10309_));
 sky130_fd_sc_hd__xnor2_1 _17802_ (.A(_10289_),
    .B(_10309_),
    .Y(_10310_));
 sky130_fd_sc_hd__and2b_1 _17803_ (.A_N(_10256_),
    .B(_10254_),
    .X(_10311_));
 sky130_fd_sc_hd__a21oi_1 _17804_ (.A1(_10239_),
    .A2(_10257_),
    .B1(_10311_),
    .Y(_10312_));
 sky130_fd_sc_hd__xnor2_1 _17805_ (.A(_10310_),
    .B(_10312_),
    .Y(_10313_));
 sky130_fd_sc_hd__xor2_1 _17806_ (.A(_10282_),
    .B(_10313_),
    .X(_10314_));
 sky130_fd_sc_hd__nor2_1 _17807_ (.A(_10258_),
    .B(_10260_),
    .Y(_10315_));
 sky130_fd_sc_hd__a21oi_1 _17808_ (.A1(_10231_),
    .A2(_10261_),
    .B1(_10315_),
    .Y(_10316_));
 sky130_fd_sc_hd__nor2_1 _17809_ (.A(_10314_),
    .B(_10316_),
    .Y(_10317_));
 sky130_fd_sc_hd__and2_1 _17810_ (.A(_10314_),
    .B(_10316_),
    .X(_10318_));
 sky130_fd_sc_hd__nor2_1 _17811_ (.A(_10317_),
    .B(_10318_),
    .Y(_10319_));
 sky130_fd_sc_hd__xnor2_1 _17812_ (.A(_10279_),
    .B(_10319_),
    .Y(_10320_));
 sky130_fd_sc_hd__nor2_1 _17813_ (.A(_10278_),
    .B(_10320_),
    .Y(_10321_));
 sky130_fd_sc_hd__a21o_1 _17814_ (.A1(_10278_),
    .A2(_10320_),
    .B1(_09292_),
    .X(_10322_));
 sky130_fd_sc_hd__o221a_1 _17815_ (.A1(net1016),
    .A2(_09266_),
    .B1(_10321_),
    .B2(_10322_),
    .C1(_09886_),
    .X(_00614_));
 sky130_fd_sc_hd__a21o_1 _17816_ (.A1(_10271_),
    .A2(_10273_),
    .B1(_10319_),
    .X(_10323_));
 sky130_fd_sc_hd__a22o_1 _17817_ (.A1(_10279_),
    .A2(_10319_),
    .B1(_10323_),
    .B2(_10278_),
    .X(_10324_));
 sky130_fd_sc_hd__or2_1 _17818_ (.A(_10310_),
    .B(_10312_),
    .X(_10325_));
 sky130_fd_sc_hd__or2b_1 _17819_ (.A(_10313_),
    .B_N(_10282_),
    .X(_10326_));
 sky130_fd_sc_hd__a21o_1 _17820_ (.A1(_10284_),
    .A2(_10288_),
    .B1(_10286_),
    .X(_10327_));
 sky130_fd_sc_hd__a21o_1 _17821_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[9] ),
    .A2(_10236_),
    .B1(_10283_),
    .X(_10328_));
 sky130_fd_sc_hd__a31o_1 _17822_ (.A1(_10040_),
    .A2(_10047_),
    .A3(_10292_),
    .B1(_10293_),
    .X(_10329_));
 sky130_fd_sc_hd__xnor2_2 _17823_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[10] ),
    .B(_10236_),
    .Y(_10330_));
 sky130_fd_sc_hd__xnor2_2 _17824_ (.A(_10329_),
    .B(_10330_),
    .Y(_10331_));
 sky130_fd_sc_hd__xnor2_2 _17825_ (.A(_10328_),
    .B(_10331_),
    .Y(_10332_));
 sky130_fd_sc_hd__or2b_1 _17826_ (.A(_10304_),
    .B_N(_10303_),
    .X(_10333_));
 sky130_fd_sc_hd__or2b_1 _17827_ (.A(_10297_),
    .B_N(_10305_),
    .X(_10334_));
 sky130_fd_sc_hd__and3_1 _17828_ (.A(\top_inst.grid_inst.data_path_wires[11][7] ),
    .B(_10052_),
    .C(_10050_),
    .X(_10335_));
 sky130_fd_sc_hd__a22o_1 _17829_ (.A1(_10037_),
    .A2(_10052_),
    .B1(_10050_),
    .B2(\top_inst.grid_inst.data_path_wires[11][7] ),
    .X(_10336_));
 sky130_fd_sc_hd__a21bo_1 _17830_ (.A1(_10038_),
    .A2(_10335_),
    .B1_N(_10336_),
    .X(_10337_));
 sky130_fd_sc_hd__xor2_1 _17831_ (.A(_10296_),
    .B(_10337_),
    .X(_10338_));
 sky130_fd_sc_hd__nand2_1 _17832_ (.A(_10035_),
    .B(_10054_),
    .Y(_10339_));
 sky130_fd_sc_hd__and4b_1 _17833_ (.A_N(\top_inst.grid_inst.data_path_wires[11][3] ),
    .B(_10059_),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[6] ),
    .D(\top_inst.grid_inst.data_path_wires[11][4] ),
    .X(_10340_));
 sky130_fd_sc_hd__o2bb2a_1 _17834_ (.A1_N(\top_inst.grid_inst.data_path_wires[11][4] ),
    .A2_N(_10056_),
    .B1(_10300_),
    .B2(\top_inst.grid_inst.data_path_wires[11][3] ),
    .X(_10341_));
 sky130_fd_sc_hd__nor2_1 _17835_ (.A(_10340_),
    .B(_10341_),
    .Y(_10342_));
 sky130_fd_sc_hd__xnor2_1 _17836_ (.A(_10339_),
    .B(_10342_),
    .Y(_10343_));
 sky130_fd_sc_hd__o21ba_1 _17837_ (.A1(_10298_),
    .A2(_10301_),
    .B1_N(_10299_),
    .X(_10344_));
 sky130_fd_sc_hd__xnor2_1 _17838_ (.A(_10343_),
    .B(_10344_),
    .Y(_10345_));
 sky130_fd_sc_hd__xnor2_1 _17839_ (.A(_10338_),
    .B(_10345_),
    .Y(_10346_));
 sky130_fd_sc_hd__a21oi_1 _17840_ (.A1(_10333_),
    .A2(_10334_),
    .B1(_10346_),
    .Y(_10347_));
 sky130_fd_sc_hd__and3_1 _17841_ (.A(_10333_),
    .B(_10334_),
    .C(_10346_),
    .X(_10348_));
 sky130_fd_sc_hd__or2_1 _17842_ (.A(_10347_),
    .B(_10348_),
    .X(_10349_));
 sky130_fd_sc_hd__xnor2_1 _17843_ (.A(_10332_),
    .B(_10349_),
    .Y(_10350_));
 sky130_fd_sc_hd__a21oi_1 _17844_ (.A1(_10289_),
    .A2(_10309_),
    .B1(_10307_),
    .Y(_10351_));
 sky130_fd_sc_hd__xnor2_1 _17845_ (.A(_10350_),
    .B(_10351_),
    .Y(_10352_));
 sky130_fd_sc_hd__xor2_1 _17846_ (.A(_10327_),
    .B(_10352_),
    .X(_10353_));
 sky130_fd_sc_hd__a21o_1 _17847_ (.A1(_10325_),
    .A2(_10326_),
    .B1(_10353_),
    .X(_10354_));
 sky130_fd_sc_hd__nand3_1 _17848_ (.A(_10325_),
    .B(_10326_),
    .C(_10353_),
    .Y(_10355_));
 sky130_fd_sc_hd__and2_1 _17849_ (.A(_10354_),
    .B(_10355_),
    .X(_10356_));
 sky130_fd_sc_hd__nand2_1 _17850_ (.A(_10317_),
    .B(_10356_),
    .Y(_10357_));
 sky130_fd_sc_hd__or2_1 _17851_ (.A(_10317_),
    .B(_10356_),
    .X(_10358_));
 sky130_fd_sc_hd__and2_1 _17852_ (.A(_10357_),
    .B(_10358_),
    .X(_10359_));
 sky130_fd_sc_hd__nand2_1 _17853_ (.A(_10324_),
    .B(_10359_),
    .Y(_10360_));
 sky130_fd_sc_hd__or2_1 _17854_ (.A(_10324_),
    .B(_10359_),
    .X(_10361_));
 sky130_fd_sc_hd__and2_1 _17855_ (.A(_10360_),
    .B(_10361_),
    .X(_10362_));
 sky130_fd_sc_hd__or2_1 _17856_ (.A(net1083),
    .B(_09494_),
    .X(_10363_));
 sky130_fd_sc_hd__o211a_1 _17857_ (.A1(_10071_),
    .A2(_10362_),
    .B1(_10363_),
    .C1(_10049_),
    .X(_00615_));
 sky130_fd_sc_hd__buf_4 _17858_ (.A(_06168_),
    .X(_10364_));
 sky130_fd_sc_hd__or2b_1 _17859_ (.A(_10330_),
    .B_N(_10329_),
    .X(_10365_));
 sky130_fd_sc_hd__a21bo_1 _17860_ (.A1(_10328_),
    .A2(_10331_),
    .B1_N(_10365_),
    .X(_10366_));
 sky130_fd_sc_hd__clkbuf_4 _17861_ (.A(_10236_),
    .X(_10367_));
 sky130_fd_sc_hd__a21o_1 _17862_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[10] ),
    .A2(_10367_),
    .B1(_10283_),
    .X(_10368_));
 sky130_fd_sc_hd__xnor2_1 _17863_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[11] ),
    .B(_10236_),
    .Y(_10369_));
 sky130_fd_sc_hd__a32o_1 _17864_ (.A1(_10040_),
    .A2(_10047_),
    .A3(_10336_),
    .B1(_10335_),
    .B2(_10038_),
    .X(_10370_));
 sky130_fd_sc_hd__and2b_1 _17865_ (.A_N(_10369_),
    .B(_10370_),
    .X(_10371_));
 sky130_fd_sc_hd__and2b_1 _17866_ (.A_N(_10370_),
    .B(_10369_),
    .X(_10372_));
 sky130_fd_sc_hd__nor2_1 _17867_ (.A(_10371_),
    .B(_10372_),
    .Y(_10373_));
 sky130_fd_sc_hd__xnor2_2 _17868_ (.A(_10368_),
    .B(_10373_),
    .Y(_10374_));
 sky130_fd_sc_hd__o21ai_1 _17869_ (.A1(_10052_),
    .A2(_10050_),
    .B1(_10040_),
    .Y(_10375_));
 sky130_fd_sc_hd__nor2_2 _17870_ (.A(_10335_),
    .B(_10375_),
    .Y(_10376_));
 sky130_fd_sc_hd__xnor2_4 _17871_ (.A(_10296_),
    .B(_10376_),
    .Y(_10377_));
 sky130_fd_sc_hd__inv_2 _17872_ (.A(\top_inst.grid_inst.data_path_wires[11][4] ),
    .Y(_10378_));
 sky130_fd_sc_hd__and4_1 _17873_ (.A(_10035_),
    .B(_10378_),
    .C(_10059_),
    .D(_10056_),
    .X(_10379_));
 sky130_fd_sc_hd__a22o_1 _17874_ (.A1(_10378_),
    .A2(_10059_),
    .B1(_10056_),
    .B2(\top_inst.grid_inst.data_path_wires[11][5] ),
    .X(_10380_));
 sky130_fd_sc_hd__and4b_1 _17875_ (.A_N(_10379_),
    .B(_10380_),
    .C(_10038_),
    .D(_10054_),
    .X(_10381_));
 sky130_fd_sc_hd__inv_2 _17876_ (.A(_10380_),
    .Y(_10382_));
 sky130_fd_sc_hd__o2bb2a_1 _17877_ (.A1_N(_10038_),
    .A2_N(_10054_),
    .B1(_10379_),
    .B2(_10382_),
    .X(_10383_));
 sky130_fd_sc_hd__nor2_1 _17878_ (.A(_10381_),
    .B(_10383_),
    .Y(_10384_));
 sky130_fd_sc_hd__o21ba_1 _17879_ (.A1(_10339_),
    .A2(_10341_),
    .B1_N(_10340_),
    .X(_10385_));
 sky130_fd_sc_hd__xnor2_1 _17880_ (.A(_10384_),
    .B(_10385_),
    .Y(_10386_));
 sky130_fd_sc_hd__xnor2_1 _17881_ (.A(_10377_),
    .B(_10386_),
    .Y(_10387_));
 sky130_fd_sc_hd__or2b_1 _17882_ (.A(_10344_),
    .B_N(_10343_),
    .X(_10388_));
 sky130_fd_sc_hd__a21bo_1 _17883_ (.A1(_10338_),
    .A2(_10345_),
    .B1_N(_10388_),
    .X(_10389_));
 sky130_fd_sc_hd__xor2_1 _17884_ (.A(_10387_),
    .B(_10389_),
    .X(_10390_));
 sky130_fd_sc_hd__xor2_1 _17885_ (.A(_10374_),
    .B(_10390_),
    .X(_10391_));
 sky130_fd_sc_hd__o21bai_1 _17886_ (.A1(_10332_),
    .A2(_10348_),
    .B1_N(_10347_),
    .Y(_10392_));
 sky130_fd_sc_hd__xnor2_1 _17887_ (.A(_10391_),
    .B(_10392_),
    .Y(_10393_));
 sky130_fd_sc_hd__xor2_1 _17888_ (.A(_10366_),
    .B(_10393_),
    .X(_10394_));
 sky130_fd_sc_hd__or2b_1 _17889_ (.A(_10352_),
    .B_N(_10327_),
    .X(_10395_));
 sky130_fd_sc_hd__o21a_1 _17890_ (.A1(_10350_),
    .A2(_10351_),
    .B1(_10395_),
    .X(_10396_));
 sky130_fd_sc_hd__or2_1 _17891_ (.A(_10394_),
    .B(_10396_),
    .X(_10397_));
 sky130_fd_sc_hd__nand2_1 _17892_ (.A(_10394_),
    .B(_10396_),
    .Y(_10398_));
 sky130_fd_sc_hd__and2_1 _17893_ (.A(_10397_),
    .B(_10398_),
    .X(_10399_));
 sky130_fd_sc_hd__xnor2_1 _17894_ (.A(_10354_),
    .B(_10399_),
    .Y(_10400_));
 sky130_fd_sc_hd__a21oi_1 _17895_ (.A1(_10357_),
    .A2(_10360_),
    .B1(_10400_),
    .Y(_10401_));
 sky130_fd_sc_hd__a31o_1 _17896_ (.A1(_10357_),
    .A2(_10360_),
    .A3(_10400_),
    .B1(_07439_),
    .X(_10402_));
 sky130_fd_sc_hd__o221a_1 _17897_ (.A1(net1038),
    .A2(_10364_),
    .B1(_10401_),
    .B2(_10402_),
    .C1(_09886_),
    .X(_00616_));
 sky130_fd_sc_hd__nand2_1 _17898_ (.A(_10354_),
    .B(_10357_),
    .Y(_10403_));
 sky130_fd_sc_hd__a32o_1 _17899_ (.A1(_10324_),
    .A2(_10359_),
    .A3(_10400_),
    .B1(_10403_),
    .B2(_10399_),
    .X(_10404_));
 sky130_fd_sc_hd__nand2_1 _17900_ (.A(_10391_),
    .B(_10392_),
    .Y(_10405_));
 sky130_fd_sc_hd__or2b_1 _17901_ (.A(_10393_),
    .B_N(_10366_),
    .X(_10406_));
 sky130_fd_sc_hd__a21o_1 _17902_ (.A1(_10368_),
    .A2(_10373_),
    .B1(_10371_),
    .X(_10407_));
 sky130_fd_sc_hd__inv_2 _17903_ (.A(_10407_),
    .Y(_10408_));
 sky130_fd_sc_hd__and2b_1 _17904_ (.A_N(_10387_),
    .B(_10389_),
    .X(_10409_));
 sky130_fd_sc_hd__o21ba_1 _17905_ (.A1(_10374_),
    .A2(_10390_),
    .B1_N(_10409_),
    .X(_10410_));
 sky130_fd_sc_hd__a21o_1 _17906_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[11] ),
    .A2(_10367_),
    .B1(_10283_),
    .X(_10411_));
 sky130_fd_sc_hd__o21ba_1 _17907_ (.A1(_10296_),
    .A2(_10375_),
    .B1_N(_10335_),
    .X(_10412_));
 sky130_fd_sc_hd__clkbuf_4 _17908_ (.A(_10412_),
    .X(_10413_));
 sky130_fd_sc_hd__xnor2_1 _17909_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[12] ),
    .B(_10236_),
    .Y(_10414_));
 sky130_fd_sc_hd__nor2_1 _17910_ (.A(_10413_),
    .B(_10414_),
    .Y(_10415_));
 sky130_fd_sc_hd__and2_1 _17911_ (.A(_10412_),
    .B(_10414_),
    .X(_10416_));
 sky130_fd_sc_hd__nor2_1 _17912_ (.A(_10415_),
    .B(_10416_),
    .Y(_10417_));
 sky130_fd_sc_hd__xnor2_1 _17913_ (.A(_10411_),
    .B(_10417_),
    .Y(_10418_));
 sky130_fd_sc_hd__nand2_1 _17914_ (.A(_10040_),
    .B(_10054_),
    .Y(_10419_));
 sky130_fd_sc_hd__nor2_1 _17915_ (.A(_10035_),
    .B(_10300_),
    .Y(_10420_));
 sky130_fd_sc_hd__and3_1 _17916_ (.A(_10037_),
    .B(_10056_),
    .C(_10420_),
    .X(_10421_));
 sky130_fd_sc_hd__a21oi_1 _17917_ (.A1(_10038_),
    .A2(_10056_),
    .B1(_10420_),
    .Y(_10422_));
 sky130_fd_sc_hd__nor3_1 _17918_ (.A(_10419_),
    .B(_10421_),
    .C(_10422_),
    .Y(_10423_));
 sky130_fd_sc_hd__o21a_1 _17919_ (.A1(_10421_),
    .A2(_10422_),
    .B1(_10419_),
    .X(_10424_));
 sky130_fd_sc_hd__nor2_1 _17920_ (.A(_10423_),
    .B(_10424_),
    .Y(_10425_));
 sky130_fd_sc_hd__nor2_1 _17921_ (.A(_10379_),
    .B(_10381_),
    .Y(_10426_));
 sky130_fd_sc_hd__xnor2_1 _17922_ (.A(_10425_),
    .B(_10426_),
    .Y(_10427_));
 sky130_fd_sc_hd__nand2_1 _17923_ (.A(_10377_),
    .B(_10427_),
    .Y(_10428_));
 sky130_fd_sc_hd__or2_1 _17924_ (.A(_10377_),
    .B(_10427_),
    .X(_10429_));
 sky130_fd_sc_hd__nand2_1 _17925_ (.A(_10428_),
    .B(_10429_),
    .Y(_10430_));
 sky130_fd_sc_hd__or3_1 _17926_ (.A(_10381_),
    .B(_10383_),
    .C(_10385_),
    .X(_10431_));
 sky130_fd_sc_hd__a21bo_1 _17927_ (.A1(_10377_),
    .A2(_10386_),
    .B1_N(_10431_),
    .X(_10432_));
 sky130_fd_sc_hd__xor2_1 _17928_ (.A(_10430_),
    .B(_10432_),
    .X(_10433_));
 sky130_fd_sc_hd__xor2_1 _17929_ (.A(_10418_),
    .B(_10433_),
    .X(_10434_));
 sky130_fd_sc_hd__or2b_1 _17930_ (.A(_10410_),
    .B_N(_10434_),
    .X(_10435_));
 sky130_fd_sc_hd__or2b_1 _17931_ (.A(_10434_),
    .B_N(_10410_),
    .X(_10436_));
 sky130_fd_sc_hd__nand2_1 _17932_ (.A(_10435_),
    .B(_10436_),
    .Y(_10437_));
 sky130_fd_sc_hd__xnor2_1 _17933_ (.A(_10408_),
    .B(_10437_),
    .Y(_10438_));
 sky130_fd_sc_hd__a21oi_1 _17934_ (.A1(_10405_),
    .A2(_10406_),
    .B1(_10438_),
    .Y(_10439_));
 sky130_fd_sc_hd__and3_1 _17935_ (.A(_10405_),
    .B(_10406_),
    .C(_10438_),
    .X(_10440_));
 sky130_fd_sc_hd__nor2_1 _17936_ (.A(_10439_),
    .B(_10440_),
    .Y(_10441_));
 sky130_fd_sc_hd__xnor2_1 _17937_ (.A(_10397_),
    .B(_10441_),
    .Y(_10442_));
 sky130_fd_sc_hd__nand2_1 _17938_ (.A(_10404_),
    .B(_10442_),
    .Y(_10443_));
 sky130_fd_sc_hd__or2_1 _17939_ (.A(_10404_),
    .B(_10442_),
    .X(_10444_));
 sky130_fd_sc_hd__and2_1 _17940_ (.A(_10443_),
    .B(_10444_),
    .X(_10445_));
 sky130_fd_sc_hd__or2_1 _17941_ (.A(net1089),
    .B(_09494_),
    .X(_10446_));
 sky130_fd_sc_hd__buf_4 _17942_ (.A(_04868_),
    .X(_10447_));
 sky130_fd_sc_hd__buf_4 _17943_ (.A(_10447_),
    .X(_10448_));
 sky130_fd_sc_hd__o211a_1 _17944_ (.A1(_10071_),
    .A2(_10445_),
    .B1(_10446_),
    .C1(_10448_),
    .X(_00617_));
 sky130_fd_sc_hd__or3_1 _17945_ (.A(_10397_),
    .B(_10439_),
    .C(_10440_),
    .X(_10449_));
 sky130_fd_sc_hd__a21o_1 _17946_ (.A1(_10405_),
    .A2(_10406_),
    .B1(_10438_),
    .X(_10450_));
 sky130_fd_sc_hd__a21o_1 _17947_ (.A1(_10411_),
    .A2(_10417_),
    .B1(_10415_),
    .X(_10451_));
 sky130_fd_sc_hd__a21o_1 _17948_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[12] ),
    .A2(_10367_),
    .B1(_10283_),
    .X(_10452_));
 sky130_fd_sc_hd__xnor2_1 _17949_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[13] ),
    .B(_10367_),
    .Y(_10453_));
 sky130_fd_sc_hd__nor2_1 _17950_ (.A(_10413_),
    .B(_10453_),
    .Y(_10454_));
 sky130_fd_sc_hd__and2_1 _17951_ (.A(_10413_),
    .B(_10453_),
    .X(_10455_));
 sky130_fd_sc_hd__nor2_1 _17952_ (.A(_10454_),
    .B(_10455_),
    .Y(_10456_));
 sky130_fd_sc_hd__xnor2_2 _17953_ (.A(_10452_),
    .B(_10456_),
    .Y(_10457_));
 sky130_fd_sc_hd__or3_1 _17954_ (.A(_10423_),
    .B(_10424_),
    .C(_10426_),
    .X(_10458_));
 sky130_fd_sc_hd__nand2_1 _17955_ (.A(\top_inst.grid_inst.data_path_wires[11][7] ),
    .B(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[6] ),
    .Y(_10459_));
 sky130_fd_sc_hd__or3_1 _17956_ (.A(_10037_),
    .B(_10300_),
    .C(_10459_),
    .X(_10460_));
 sky130_fd_sc_hd__o21ai_1 _17957_ (.A1(_10037_),
    .A2(_10300_),
    .B1(_10459_),
    .Y(_10461_));
 sky130_fd_sc_hd__and2_1 _17958_ (.A(_10460_),
    .B(_10461_),
    .X(_10462_));
 sky130_fd_sc_hd__xnor2_1 _17959_ (.A(_10419_),
    .B(_10462_),
    .Y(_10463_));
 sky130_fd_sc_hd__o21ai_1 _17960_ (.A1(_10421_),
    .A2(_10423_),
    .B1(_10463_),
    .Y(_10464_));
 sky130_fd_sc_hd__or3_1 _17961_ (.A(_10421_),
    .B(_10423_),
    .C(_10463_),
    .X(_10465_));
 sky130_fd_sc_hd__and2_1 _17962_ (.A(_10464_),
    .B(_10465_),
    .X(_10466_));
 sky130_fd_sc_hd__nand2_1 _17963_ (.A(_10377_),
    .B(_10466_),
    .Y(_10467_));
 sky130_fd_sc_hd__or2_1 _17964_ (.A(_10377_),
    .B(_10466_),
    .X(_10468_));
 sky130_fd_sc_hd__nand2_1 _17965_ (.A(_10467_),
    .B(_10468_),
    .Y(_10469_));
 sky130_fd_sc_hd__a21o_1 _17966_ (.A1(_10458_),
    .A2(_10428_),
    .B1(_10469_),
    .X(_10470_));
 sky130_fd_sc_hd__nand3_1 _17967_ (.A(_10458_),
    .B(_10428_),
    .C(_10469_),
    .Y(_10471_));
 sky130_fd_sc_hd__nand2_1 _17968_ (.A(_10470_),
    .B(_10471_),
    .Y(_10472_));
 sky130_fd_sc_hd__xor2_2 _17969_ (.A(_10457_),
    .B(_10472_),
    .X(_10473_));
 sky130_fd_sc_hd__or2b_1 _17970_ (.A(_10430_),
    .B_N(_10432_),
    .X(_10474_));
 sky130_fd_sc_hd__o21a_1 _17971_ (.A1(_10418_),
    .A2(_10433_),
    .B1(_10474_),
    .X(_10475_));
 sky130_fd_sc_hd__xor2_1 _17972_ (.A(_10473_),
    .B(_10475_),
    .X(_10476_));
 sky130_fd_sc_hd__xor2_1 _17973_ (.A(_10451_),
    .B(_10476_),
    .X(_10477_));
 sky130_fd_sc_hd__o21a_1 _17974_ (.A1(_10408_),
    .A2(_10437_),
    .B1(_10435_),
    .X(_10478_));
 sky130_fd_sc_hd__or2_1 _17975_ (.A(_10477_),
    .B(_10478_),
    .X(_10479_));
 sky130_fd_sc_hd__nand2_1 _17976_ (.A(_10477_),
    .B(_10478_),
    .Y(_10480_));
 sky130_fd_sc_hd__and2_1 _17977_ (.A(_10479_),
    .B(_10480_),
    .X(_10481_));
 sky130_fd_sc_hd__xnor2_1 _17978_ (.A(_10450_),
    .B(_10481_),
    .Y(_10482_));
 sky130_fd_sc_hd__a21oi_1 _17979_ (.A1(_10449_),
    .A2(_10443_),
    .B1(_10482_),
    .Y(_10483_));
 sky130_fd_sc_hd__a31o_1 _17980_ (.A1(_10449_),
    .A2(_10443_),
    .A3(_10482_),
    .B1(_07439_),
    .X(_10484_));
 sky130_fd_sc_hd__o221a_1 _17981_ (.A1(net1011),
    .A2(_10364_),
    .B1(_10483_),
    .B2(_10484_),
    .C1(_09886_),
    .X(_00618_));
 sky130_fd_sc_hd__nand2_1 _17982_ (.A(_10450_),
    .B(_10449_),
    .Y(_10485_));
 sky130_fd_sc_hd__a32o_1 _17983_ (.A1(_10404_),
    .A2(_10442_),
    .A3(_10482_),
    .B1(_10485_),
    .B2(_10481_),
    .X(_10486_));
 sky130_fd_sc_hd__a21o_1 _17984_ (.A1(_10452_),
    .A2(_10456_),
    .B1(_10454_),
    .X(_10487_));
 sky130_fd_sc_hd__inv_2 _17985_ (.A(_10487_),
    .Y(_10488_));
 sky130_fd_sc_hd__o21a_1 _17986_ (.A1(_10457_),
    .A2(_10472_),
    .B1(_10470_),
    .X(_10489_));
 sky130_fd_sc_hd__a21o_1 _17987_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[13] ),
    .A2(_10367_),
    .B1(_10283_),
    .X(_10490_));
 sky130_fd_sc_hd__and2_1 _17988_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[14] ),
    .B(_10367_),
    .X(_10491_));
 sky130_fd_sc_hd__nor2_1 _17989_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[14] ),
    .B(_10367_),
    .Y(_10492_));
 sky130_fd_sc_hd__or2_1 _17990_ (.A(_10491_),
    .B(_10492_),
    .X(_10493_));
 sky130_fd_sc_hd__xor2_1 _17991_ (.A(_10413_),
    .B(_10493_),
    .X(_10494_));
 sky130_fd_sc_hd__nand2_1 _17992_ (.A(_10490_),
    .B(_10494_),
    .Y(_10495_));
 sky130_fd_sc_hd__or2_1 _17993_ (.A(_10490_),
    .B(_10494_),
    .X(_10496_));
 sky130_fd_sc_hd__nand2_1 _17994_ (.A(_10495_),
    .B(_10496_),
    .Y(_10497_));
 sky130_fd_sc_hd__o211a_1 _17995_ (.A1(_10040_),
    .A2(_10300_),
    .B1(_10419_),
    .C1(_10459_),
    .X(_10498_));
 sky130_fd_sc_hd__and2_1 _17996_ (.A(_10040_),
    .B(_10054_),
    .X(_10499_));
 sky130_fd_sc_hd__nand2_1 _17997_ (.A(_10499_),
    .B(_10462_),
    .Y(_10500_));
 sky130_fd_sc_hd__a22oi_2 _17998_ (.A1(_10056_),
    .A2(_10499_),
    .B1(_10460_),
    .B2(_10500_),
    .Y(_10501_));
 sky130_fd_sc_hd__nor2_1 _17999_ (.A(_10498_),
    .B(_10501_),
    .Y(_10502_));
 sky130_fd_sc_hd__xnor2_1 _18000_ (.A(_10377_),
    .B(_10502_),
    .Y(_10503_));
 sky130_fd_sc_hd__a21oi_1 _18001_ (.A1(_10464_),
    .A2(_10467_),
    .B1(_10503_),
    .Y(_10504_));
 sky130_fd_sc_hd__and3_1 _18002_ (.A(_10464_),
    .B(_10467_),
    .C(_10503_),
    .X(_10505_));
 sky130_fd_sc_hd__nor2_1 _18003_ (.A(_10504_),
    .B(_10505_),
    .Y(_10506_));
 sky130_fd_sc_hd__xnor2_1 _18004_ (.A(_10497_),
    .B(_10506_),
    .Y(_10507_));
 sky130_fd_sc_hd__or2b_1 _18005_ (.A(_10489_),
    .B_N(_10507_),
    .X(_10508_));
 sky130_fd_sc_hd__or2b_1 _18006_ (.A(_10507_),
    .B_N(_10489_),
    .X(_10509_));
 sky130_fd_sc_hd__nand2_1 _18007_ (.A(_10508_),
    .B(_10509_),
    .Y(_10510_));
 sky130_fd_sc_hd__xnor2_2 _18008_ (.A(_10488_),
    .B(_10510_),
    .Y(_10511_));
 sky130_fd_sc_hd__inv_2 _18009_ (.A(_10475_),
    .Y(_10512_));
 sky130_fd_sc_hd__and2b_1 _18010_ (.A_N(_10476_),
    .B(_10451_),
    .X(_10513_));
 sky130_fd_sc_hd__a21oi_2 _18011_ (.A1(_10473_),
    .A2(_10512_),
    .B1(_10513_),
    .Y(_10514_));
 sky130_fd_sc_hd__xor2_2 _18012_ (.A(_10511_),
    .B(_10514_),
    .X(_10515_));
 sky130_fd_sc_hd__xnor2_2 _18013_ (.A(_10479_),
    .B(_10515_),
    .Y(_10516_));
 sky130_fd_sc_hd__xor2_1 _18014_ (.A(_10486_),
    .B(_10516_),
    .X(_10517_));
 sky130_fd_sc_hd__or2_1 _18015_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[14] ),
    .B(_09494_),
    .X(_10518_));
 sky130_fd_sc_hd__o211a_1 _18016_ (.A1(_10071_),
    .A2(_10517_),
    .B1(_10518_),
    .C1(_10448_),
    .X(_00619_));
 sky130_fd_sc_hd__or2b_1 _18017_ (.A(_10479_),
    .B_N(_10515_),
    .X(_10519_));
 sky130_fd_sc_hd__a21boi_1 _18018_ (.A1(_10486_),
    .A2(_10516_),
    .B1_N(_10519_),
    .Y(_10520_));
 sky130_fd_sc_hd__or2_1 _18019_ (.A(_10511_),
    .B(_10514_),
    .X(_10521_));
 sky130_fd_sc_hd__o21ai_1 _18020_ (.A1(_10413_),
    .A2(_10493_),
    .B1(_10495_),
    .Y(_10522_));
 sky130_fd_sc_hd__nor2_1 _18021_ (.A(_10377_),
    .B(_10502_),
    .Y(_10523_));
 sky130_fd_sc_hd__xnor2_1 _18022_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[15] ),
    .B(_10367_),
    .Y(_10524_));
 sky130_fd_sc_hd__nor2_1 _18023_ (.A(_10413_),
    .B(_10524_),
    .Y(_10525_));
 sky130_fd_sc_hd__and2_1 _18024_ (.A(_10413_),
    .B(_10524_),
    .X(_10526_));
 sky130_fd_sc_hd__nor2_1 _18025_ (.A(_10525_),
    .B(_10526_),
    .Y(_10527_));
 sky130_fd_sc_hd__o21a_1 _18026_ (.A1(_10283_),
    .A2(_10491_),
    .B1(_10527_),
    .X(_10528_));
 sky130_fd_sc_hd__nor3_1 _18027_ (.A(_10283_),
    .B(_10491_),
    .C(_10527_),
    .Y(_10529_));
 sky130_fd_sc_hd__or2_1 _18028_ (.A(_10528_),
    .B(_10529_),
    .X(_10530_));
 sky130_fd_sc_hd__xor2_1 _18029_ (.A(_10523_),
    .B(_10530_),
    .X(_10531_));
 sky130_fd_sc_hd__a31o_1 _18030_ (.A1(_10495_),
    .A2(_10496_),
    .A3(_10506_),
    .B1(_10504_),
    .X(_10532_));
 sky130_fd_sc_hd__xnor2_1 _18031_ (.A(_10531_),
    .B(_10532_),
    .Y(_10533_));
 sky130_fd_sc_hd__xor2_1 _18032_ (.A(_10522_),
    .B(_10533_),
    .X(_10534_));
 sky130_fd_sc_hd__o21a_1 _18033_ (.A1(_10488_),
    .A2(_10510_),
    .B1(_10508_),
    .X(_10535_));
 sky130_fd_sc_hd__or2_1 _18034_ (.A(_10534_),
    .B(_10535_),
    .X(_10536_));
 sky130_fd_sc_hd__nand2_1 _18035_ (.A(_10534_),
    .B(_10535_),
    .Y(_10537_));
 sky130_fd_sc_hd__and2_1 _18036_ (.A(_10536_),
    .B(_10537_),
    .X(_10538_));
 sky130_fd_sc_hd__xnor2_1 _18037_ (.A(_10521_),
    .B(_10538_),
    .Y(_10539_));
 sky130_fd_sc_hd__nor2_1 _18038_ (.A(_10520_),
    .B(_10539_),
    .Y(_10540_));
 sky130_fd_sc_hd__clkbuf_4 _18039_ (.A(_05309_),
    .X(_10541_));
 sky130_fd_sc_hd__a2111o_1 _18040_ (.A1(_10520_),
    .A2(_10539_),
    .B1(_10540_),
    .C1(_10541_),
    .D1(_04861_),
    .X(_10542_));
 sky130_fd_sc_hd__o211a_1 _18041_ (.A1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[15] ),
    .A2(_08183_),
    .B1(_10542_),
    .C1(_10448_),
    .X(_00620_));
 sky130_fd_sc_hd__nand2_1 _18042_ (.A(_10521_),
    .B(_10519_),
    .Y(_10543_));
 sky130_fd_sc_hd__a32o_1 _18043_ (.A1(_10486_),
    .A2(_10516_),
    .A3(_10539_),
    .B1(_10543_),
    .B2(_10538_),
    .X(_10544_));
 sky130_fd_sc_hd__inv_2 _18044_ (.A(_10377_),
    .Y(_10545_));
 sky130_fd_sc_hd__o2bb2a_1 _18045_ (.A1_N(_10545_),
    .A2_N(_10501_),
    .B1(_10523_),
    .B2(_10530_),
    .X(_10546_));
 sky130_fd_sc_hd__nand2_1 _18046_ (.A(_10545_),
    .B(_10498_),
    .Y(_10547_));
 sky130_fd_sc_hd__a21o_1 _18047_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[15] ),
    .A2(_10367_),
    .B1(_10283_),
    .X(_10548_));
 sky130_fd_sc_hd__xnor2_1 _18048_ (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[16] ),
    .B(_10367_),
    .Y(_10549_));
 sky130_fd_sc_hd__xor2_1 _18049_ (.A(_10413_),
    .B(_10549_),
    .X(_10550_));
 sky130_fd_sc_hd__xnor2_1 _18050_ (.A(_10548_),
    .B(_10550_),
    .Y(_10551_));
 sky130_fd_sc_hd__xor2_1 _18051_ (.A(_10547_),
    .B(_10551_),
    .X(_10552_));
 sky130_fd_sc_hd__xor2_1 _18052_ (.A(_10546_),
    .B(_10552_),
    .X(_10553_));
 sky130_fd_sc_hd__o21ai_1 _18053_ (.A1(_10525_),
    .A2(_10528_),
    .B1(_10553_),
    .Y(_10554_));
 sky130_fd_sc_hd__or3_1 _18054_ (.A(_10525_),
    .B(_10528_),
    .C(_10553_),
    .X(_10555_));
 sky130_fd_sc_hd__nand2_1 _18055_ (.A(_10554_),
    .B(_10555_),
    .Y(_10556_));
 sky130_fd_sc_hd__and2b_1 _18056_ (.A_N(_10533_),
    .B(_10522_),
    .X(_10557_));
 sky130_fd_sc_hd__a21oi_1 _18057_ (.A1(_10531_),
    .A2(_10532_),
    .B1(_10557_),
    .Y(_10558_));
 sky130_fd_sc_hd__xor2_1 _18058_ (.A(_10556_),
    .B(_10558_),
    .X(_10559_));
 sky130_fd_sc_hd__xnor2_1 _18059_ (.A(_10536_),
    .B(_10559_),
    .Y(_10560_));
 sky130_fd_sc_hd__xor2_1 _18060_ (.A(_10544_),
    .B(_10560_),
    .X(_10561_));
 sky130_fd_sc_hd__or2_1 _18061_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[16] ),
    .B(_09494_),
    .X(_10562_));
 sky130_fd_sc_hd__o211a_1 _18062_ (.A1(_10071_),
    .A2(_10561_),
    .B1(_10562_),
    .C1(_10448_),
    .X(_00621_));
 sky130_fd_sc_hd__clkbuf_4 _18063_ (.A(_05313_),
    .X(_10563_));
 sky130_fd_sc_hd__nor2_1 _18064_ (.A(_10556_),
    .B(_10558_),
    .Y(_10564_));
 sky130_fd_sc_hd__o21a_1 _18065_ (.A1(_10546_),
    .A2(_10552_),
    .B1(_10554_),
    .X(_10565_));
 sky130_fd_sc_hd__a21o_1 _18066_ (.A1(_10413_),
    .A2(_10549_),
    .B1(_10548_),
    .X(_10566_));
 sky130_fd_sc_hd__o21a_1 _18067_ (.A1(_10413_),
    .A2(_10549_),
    .B1(_10566_),
    .X(_10567_));
 sky130_fd_sc_hd__nand2_1 _18068_ (.A(_10547_),
    .B(_10551_),
    .Y(_10568_));
 sky130_fd_sc_hd__o21ba_1 _18069_ (.A1(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[16] ),
    .A2(_10283_),
    .B1_N(_10234_),
    .X(_10569_));
 sky130_fd_sc_hd__xnor2_1 _18070_ (.A(_10568_),
    .B(_10569_),
    .Y(_10570_));
 sky130_fd_sc_hd__xnor2_1 _18071_ (.A(_10567_),
    .B(_10570_),
    .Y(_10571_));
 sky130_fd_sc_hd__xnor2_1 _18072_ (.A(_10565_),
    .B(_10571_),
    .Y(_10572_));
 sky130_fd_sc_hd__xnor2_1 _18073_ (.A(_10564_),
    .B(_10572_),
    .Y(_10573_));
 sky130_fd_sc_hd__and2b_1 _18074_ (.A_N(_10536_),
    .B(_10559_),
    .X(_10574_));
 sky130_fd_sc_hd__a211o_1 _18075_ (.A1(_10544_),
    .A2(_10560_),
    .B1(_10573_),
    .C1(_10574_),
    .X(_10575_));
 sky130_fd_sc_hd__a21oi_4 _18076_ (.A1(_05787_),
    .A2(_10575_),
    .B1(_04867_),
    .Y(_10576_));
 sky130_fd_sc_hd__o21a_1 _18077_ (.A1(net946),
    .A2(_10563_),
    .B1(_10576_),
    .X(_00622_));
 sky130_fd_sc_hd__o21a_1 _18078_ (.A1(net956),
    .A2(_10563_),
    .B1(_10576_),
    .X(_00623_));
 sky130_fd_sc_hd__o21a_1 _18079_ (.A1(net928),
    .A2(_10563_),
    .B1(_10576_),
    .X(_00624_));
 sky130_fd_sc_hd__o21a_1 _18080_ (.A1(net1002),
    .A2(_10563_),
    .B1(_10576_),
    .X(_00625_));
 sky130_fd_sc_hd__o21a_1 _18081_ (.A1(net961),
    .A2(_10563_),
    .B1(_10576_),
    .X(_00626_));
 sky130_fd_sc_hd__o21a_1 _18082_ (.A1(net975),
    .A2(_10563_),
    .B1(_10576_),
    .X(_00627_));
 sky130_fd_sc_hd__o21a_1 _18083_ (.A1(net639),
    .A2(_10563_),
    .B1(_10576_),
    .X(_00628_));
 sky130_fd_sc_hd__o21a_1 _18084_ (.A1(net1076),
    .A2(_10563_),
    .B1(_10576_),
    .X(_00629_));
 sky130_fd_sc_hd__o21a_1 _18085_ (.A1(net859),
    .A2(_10563_),
    .B1(_10576_),
    .X(_00630_));
 sky130_fd_sc_hd__o21a_1 _18086_ (.A1(net646),
    .A2(_10563_),
    .B1(_10576_),
    .X(_00631_));
 sky130_fd_sc_hd__clkbuf_4 _18087_ (.A(\top_inst.grid_inst.data_path_wires[12][0] ),
    .X(_10577_));
 sky130_fd_sc_hd__or2_1 _18088_ (.A(_10577_),
    .B(_08674_),
    .X(_10578_));
 sky130_fd_sc_hd__o211a_1 _18089_ (.A1(_10022_),
    .A2(_08663_),
    .B1(_10578_),
    .C1(_10448_),
    .X(_00632_));
 sky130_fd_sc_hd__inv_2 _18090_ (.A(\top_inst.grid_inst.data_path_wires[12][1] ),
    .Y(_10579_));
 sky130_fd_sc_hd__nand2_1 _18091_ (.A(_10579_),
    .B(_04859_),
    .Y(_10580_));
 sky130_fd_sc_hd__o211a_1 _18092_ (.A1(_10025_),
    .A2(_08663_),
    .B1(_10580_),
    .C1(_10448_),
    .X(_00633_));
 sky130_fd_sc_hd__clkbuf_4 _18093_ (.A(\top_inst.grid_inst.data_path_wires[12][2] ),
    .X(_10581_));
 sky130_fd_sc_hd__or2_1 _18094_ (.A(_10581_),
    .B(_08674_),
    .X(_10582_));
 sky130_fd_sc_hd__o211a_1 _18095_ (.A1(_10027_),
    .A2(_08663_),
    .B1(_10582_),
    .C1(_10448_),
    .X(_00634_));
 sky130_fd_sc_hd__buf_4 _18096_ (.A(_04858_),
    .X(_10583_));
 sky130_fd_sc_hd__clkbuf_4 _18097_ (.A(_10583_),
    .X(_10584_));
 sky130_fd_sc_hd__clkbuf_4 _18098_ (.A(\top_inst.grid_inst.data_path_wires[12][3] ),
    .X(_10585_));
 sky130_fd_sc_hd__or2_1 _18099_ (.A(_10585_),
    .B(_08674_),
    .X(_10586_));
 sky130_fd_sc_hd__o211a_1 _18100_ (.A1(_10029_),
    .A2(_10584_),
    .B1(_10586_),
    .C1(_10448_),
    .X(_00635_));
 sky130_fd_sc_hd__inv_2 _18101_ (.A(\top_inst.grid_inst.data_path_wires[12][4] ),
    .Y(_10587_));
 sky130_fd_sc_hd__nand2_1 _18102_ (.A(_10587_),
    .B(_04859_),
    .Y(_10588_));
 sky130_fd_sc_hd__o211a_1 _18103_ (.A1(_10032_),
    .A2(_10584_),
    .B1(_10588_),
    .C1(_10448_),
    .X(_00636_));
 sky130_fd_sc_hd__clkbuf_4 _18104_ (.A(\top_inst.grid_inst.data_path_wires[12][5] ),
    .X(_10589_));
 sky130_fd_sc_hd__or2_1 _18105_ (.A(_10589_),
    .B(_08674_),
    .X(_10590_));
 sky130_fd_sc_hd__o211a_1 _18106_ (.A1(_10035_),
    .A2(_10584_),
    .B1(_10590_),
    .C1(_10448_),
    .X(_00637_));
 sky130_fd_sc_hd__buf_2 _18107_ (.A(\top_inst.grid_inst.data_path_wires[12][6] ),
    .X(_10591_));
 sky130_fd_sc_hd__clkbuf_4 _18108_ (.A(_10591_),
    .X(_10592_));
 sky130_fd_sc_hd__or2_1 _18109_ (.A(_10592_),
    .B(_08674_),
    .X(_10593_));
 sky130_fd_sc_hd__clkbuf_4 _18110_ (.A(_10447_),
    .X(_10594_));
 sky130_fd_sc_hd__o211a_1 _18111_ (.A1(_10038_),
    .A2(_10584_),
    .B1(_10593_),
    .C1(_10594_),
    .X(_00638_));
 sky130_fd_sc_hd__clkbuf_4 _18112_ (.A(\top_inst.grid_inst.data_path_wires[12][7] ),
    .X(_10595_));
 sky130_fd_sc_hd__or2_1 _18113_ (.A(_10595_),
    .B(_08674_),
    .X(_10596_));
 sky130_fd_sc_hd__o211a_1 _18114_ (.A1(_10040_),
    .A2(_10584_),
    .B1(_10596_),
    .C1(_10594_),
    .X(_00639_));
 sky130_fd_sc_hd__clkbuf_4 _18115_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[0] ),
    .X(_10597_));
 sky130_fd_sc_hd__or2_1 _18116_ (.A(_10597_),
    .B(_10057_),
    .X(_10598_));
 sky130_fd_sc_hd__o211a_1 _18117_ (.A1(_10577_),
    .A2(_10046_),
    .B1(_10598_),
    .C1(_10594_),
    .X(_00640_));
 sky130_fd_sc_hd__clkbuf_4 _18118_ (.A(\top_inst.grid_inst.data_path_wires[12][1] ),
    .X(_10599_));
 sky130_fd_sc_hd__clkbuf_4 _18119_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[1] ),
    .X(_10600_));
 sky130_fd_sc_hd__or2_1 _18120_ (.A(_10600_),
    .B(_10057_),
    .X(_10601_));
 sky130_fd_sc_hd__o211a_1 _18121_ (.A1(_10599_),
    .A2(_10046_),
    .B1(_10601_),
    .C1(_10594_),
    .X(_00641_));
 sky130_fd_sc_hd__buf_4 _18122_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[2] ),
    .X(_10602_));
 sky130_fd_sc_hd__or2_1 _18123_ (.A(_10602_),
    .B(_10057_),
    .X(_10603_));
 sky130_fd_sc_hd__o211a_1 _18124_ (.A1(_10581_),
    .A2(_10046_),
    .B1(_10603_),
    .C1(_10594_),
    .X(_00642_));
 sky130_fd_sc_hd__clkbuf_4 _18125_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[3] ),
    .X(_10604_));
 sky130_fd_sc_hd__or2_1 _18126_ (.A(_10604_),
    .B(_10057_),
    .X(_10605_));
 sky130_fd_sc_hd__o211a_1 _18127_ (.A1(_10585_),
    .A2(_10046_),
    .B1(_10605_),
    .C1(_10594_),
    .X(_00643_));
 sky130_fd_sc_hd__clkbuf_4 _18128_ (.A(\top_inst.grid_inst.data_path_wires[12][4] ),
    .X(_10606_));
 sky130_fd_sc_hd__clkbuf_4 _18129_ (.A(_05755_),
    .X(_10607_));
 sky130_fd_sc_hd__clkbuf_4 _18130_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[4] ),
    .X(_10608_));
 sky130_fd_sc_hd__or2_1 _18131_ (.A(_10608_),
    .B(_10057_),
    .X(_10609_));
 sky130_fd_sc_hd__o211a_1 _18132_ (.A1(_10606_),
    .A2(_10607_),
    .B1(_10609_),
    .C1(_10594_),
    .X(_00644_));
 sky130_fd_sc_hd__clkbuf_4 _18133_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[5] ),
    .X(_10610_));
 sky130_fd_sc_hd__or2_1 _18134_ (.A(_10610_),
    .B(_10057_),
    .X(_10611_));
 sky130_fd_sc_hd__o211a_1 _18135_ (.A1(_10589_),
    .A2(_10607_),
    .B1(_10611_),
    .C1(_10594_),
    .X(_00645_));
 sky130_fd_sc_hd__buf_2 _18136_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[6] ),
    .X(_10612_));
 sky130_fd_sc_hd__or2_1 _18137_ (.A(_10612_),
    .B(_10057_),
    .X(_10613_));
 sky130_fd_sc_hd__o211a_1 _18138_ (.A1(_10592_),
    .A2(_10607_),
    .B1(_10613_),
    .C1(_10594_),
    .X(_00646_));
 sky130_fd_sc_hd__clkbuf_4 _18139_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[7] ),
    .X(_10614_));
 sky130_fd_sc_hd__or2_1 _18140_ (.A(_10614_),
    .B(_10057_),
    .X(_10615_));
 sky130_fd_sc_hd__o211a_1 _18141_ (.A1(_10595_),
    .A2(_10607_),
    .B1(_10615_),
    .C1(_10594_),
    .X(_00647_));
 sky130_fd_sc_hd__buf_4 _18142_ (.A(_05787_),
    .X(_10616_));
 sky130_fd_sc_hd__and3_1 _18143_ (.A(_10577_),
    .B(_10597_),
    .C(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[0] ),
    .X(_10617_));
 sky130_fd_sc_hd__a21oi_1 _18144_ (.A1(_10577_),
    .A2(_10597_),
    .B1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[0] ),
    .Y(_10618_));
 sky130_fd_sc_hd__o21ai_1 _18145_ (.A1(_10617_),
    .A2(_10618_),
    .B1(_08181_),
    .Y(_10619_));
 sky130_fd_sc_hd__clkbuf_4 _18146_ (.A(_10447_),
    .X(_10620_));
 sky130_fd_sc_hd__o211a_1 _18147_ (.A1(net996),
    .A2(_10616_),
    .B1(_10619_),
    .C1(_10620_),
    .X(_00648_));
 sky130_fd_sc_hd__a22o_1 _18148_ (.A1(\top_inst.grid_inst.data_path_wires[12][0] ),
    .A2(_10600_),
    .B1(_10597_),
    .B2(_10599_),
    .X(_10621_));
 sky130_fd_sc_hd__nand4_2 _18149_ (.A(_10599_),
    .B(_10577_),
    .C(_10600_),
    .D(_10597_),
    .Y(_10622_));
 sky130_fd_sc_hd__nand3_1 _18150_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[1] ),
    .B(_10621_),
    .C(_10622_),
    .Y(_10623_));
 sky130_fd_sc_hd__a21o_1 _18151_ (.A1(_10621_),
    .A2(_10622_),
    .B1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[1] ),
    .X(_10624_));
 sky130_fd_sc_hd__a21o_1 _18152_ (.A1(_10623_),
    .A2(_10624_),
    .B1(_10617_),
    .X(_10625_));
 sky130_fd_sc_hd__nand3_2 _18153_ (.A(_10617_),
    .B(_10623_),
    .C(_10624_),
    .Y(_10626_));
 sky130_fd_sc_hd__a21o_1 _18154_ (.A1(_10625_),
    .A2(_10626_),
    .B1(_06682_),
    .X(_10627_));
 sky130_fd_sc_hd__o211a_1 _18155_ (.A1(net935),
    .A2(_10616_),
    .B1(_10627_),
    .C1(_10620_),
    .X(_00649_));
 sky130_fd_sc_hd__nand2_1 _18156_ (.A(_10577_),
    .B(_10602_),
    .Y(_10628_));
 sky130_fd_sc_hd__a22o_1 _18157_ (.A1(_10599_),
    .A2(_10600_),
    .B1(_10597_),
    .B2(_10581_),
    .X(_10629_));
 sky130_fd_sc_hd__nand4_1 _18158_ (.A(_10581_),
    .B(_10599_),
    .C(_10600_),
    .D(_10597_),
    .Y(_10630_));
 sky130_fd_sc_hd__nand2_1 _18159_ (.A(_10629_),
    .B(_10630_),
    .Y(_10631_));
 sky130_fd_sc_hd__xor2_1 _18160_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[2] ),
    .B(_10631_),
    .X(_10632_));
 sky130_fd_sc_hd__nand2_1 _18161_ (.A(_10622_),
    .B(_10623_),
    .Y(_10633_));
 sky130_fd_sc_hd__xor2_1 _18162_ (.A(_10632_),
    .B(_10633_),
    .X(_10634_));
 sky130_fd_sc_hd__or2_1 _18163_ (.A(_10628_),
    .B(_10634_),
    .X(_10635_));
 sky130_fd_sc_hd__nand2_1 _18164_ (.A(_10628_),
    .B(_10634_),
    .Y(_10636_));
 sky130_fd_sc_hd__and2_1 _18165_ (.A(_10635_),
    .B(_10636_),
    .X(_10637_));
 sky130_fd_sc_hd__xnor2_1 _18166_ (.A(_10626_),
    .B(_10637_),
    .Y(_10638_));
 sky130_fd_sc_hd__clkbuf_4 _18167_ (.A(_06701_),
    .X(_10639_));
 sky130_fd_sc_hd__or2_1 _18168_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[2] ),
    .B(_10639_),
    .X(_10640_));
 sky130_fd_sc_hd__o211a_1 _18169_ (.A1(_10071_),
    .A2(_10638_),
    .B1(_10640_),
    .C1(_10620_),
    .X(_00650_));
 sky130_fd_sc_hd__buf_2 _18170_ (.A(_04873_),
    .X(_10641_));
 sky130_fd_sc_hd__or2b_1 _18171_ (.A(_10626_),
    .B_N(_10637_),
    .X(_10642_));
 sky130_fd_sc_hd__or2b_1 _18172_ (.A(_10632_),
    .B_N(_10633_),
    .X(_10643_));
 sky130_fd_sc_hd__a22o_1 _18173_ (.A1(_10577_),
    .A2(_10604_),
    .B1(_10602_),
    .B2(_10599_),
    .X(_10644_));
 sky130_fd_sc_hd__and3_1 _18174_ (.A(\top_inst.grid_inst.data_path_wires[12][1] ),
    .B(\top_inst.grid_inst.data_path_wires[12][0] ),
    .C(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[3] ),
    .X(_10645_));
 sky130_fd_sc_hd__nand2_2 _18175_ (.A(_10602_),
    .B(_10645_),
    .Y(_10646_));
 sky130_fd_sc_hd__nand2_1 _18176_ (.A(_10644_),
    .B(_10646_),
    .Y(_10647_));
 sky130_fd_sc_hd__a22o_1 _18177_ (.A1(_10581_),
    .A2(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[0] ),
    .B2(_10585_),
    .X(_10648_));
 sky130_fd_sc_hd__nand4_1 _18178_ (.A(_10585_),
    .B(_10581_),
    .C(_10600_),
    .D(_10597_),
    .Y(_10649_));
 sky130_fd_sc_hd__and3_1 _18179_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[3] ),
    .B(_10648_),
    .C(_10649_),
    .X(_10650_));
 sky130_fd_sc_hd__a21oi_1 _18180_ (.A1(_10648_),
    .A2(_10649_),
    .B1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[3] ),
    .Y(_10651_));
 sky130_fd_sc_hd__or2_1 _18181_ (.A(_10650_),
    .B(_10651_),
    .X(_10652_));
 sky130_fd_sc_hd__a21boi_2 _18182_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[2] ),
    .A2(_10629_),
    .B1_N(_10630_),
    .Y(_10653_));
 sky130_fd_sc_hd__xnor2_1 _18183_ (.A(_10652_),
    .B(_10653_),
    .Y(_10654_));
 sky130_fd_sc_hd__xnor2_1 _18184_ (.A(_10647_),
    .B(_10654_),
    .Y(_10655_));
 sky130_fd_sc_hd__a21o_1 _18185_ (.A1(_10643_),
    .A2(_10635_),
    .B1(_10655_),
    .X(_10656_));
 sky130_fd_sc_hd__inv_2 _18186_ (.A(_10656_),
    .Y(_10657_));
 sky130_fd_sc_hd__and3_1 _18187_ (.A(_10643_),
    .B(_10635_),
    .C(_10655_),
    .X(_10658_));
 sky130_fd_sc_hd__or3_1 _18188_ (.A(_10642_),
    .B(_10657_),
    .C(_10658_),
    .X(_10659_));
 sky130_fd_sc_hd__o21ai_1 _18189_ (.A1(_10657_),
    .A2(_10658_),
    .B1(_10642_),
    .Y(_10660_));
 sky130_fd_sc_hd__and2_1 _18190_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[3] ),
    .B(_05730_),
    .X(_10661_));
 sky130_fd_sc_hd__a31o_1 _18191_ (.A1(_05887_),
    .A2(_10659_),
    .A3(_10660_),
    .B1(_10661_),
    .X(_10662_));
 sky130_fd_sc_hd__and2_1 _18192_ (.A(_10641_),
    .B(_10662_),
    .X(_10663_));
 sky130_fd_sc_hd__clkbuf_1 _18193_ (.A(_10663_),
    .X(_00651_));
 sky130_fd_sc_hd__a22o_1 _18194_ (.A1(\top_inst.grid_inst.data_path_wires[12][3] ),
    .A2(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[12][4] ),
    .X(_10664_));
 sky130_fd_sc_hd__nand4_1 _18195_ (.A(_10606_),
    .B(_10585_),
    .C(_10600_),
    .D(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[0] ),
    .Y(_10665_));
 sky130_fd_sc_hd__nand2_1 _18196_ (.A(_10664_),
    .B(_10665_),
    .Y(_10666_));
 sky130_fd_sc_hd__xor2_2 _18197_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[4] ),
    .B(_10666_),
    .X(_10667_));
 sky130_fd_sc_hd__xor2_2 _18198_ (.A(_10646_),
    .B(_10667_),
    .X(_10668_));
 sky130_fd_sc_hd__a21bo_1 _18199_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[3] ),
    .A2(_10648_),
    .B1_N(_10649_),
    .X(_10669_));
 sky130_fd_sc_hd__xnor2_2 _18200_ (.A(_10668_),
    .B(_10669_),
    .Y(_10670_));
 sky130_fd_sc_hd__nand2_1 _18201_ (.A(_10581_),
    .B(_10602_),
    .Y(_10671_));
 sky130_fd_sc_hd__a22o_1 _18202_ (.A1(\top_inst.grid_inst.data_path_wires[12][0] ),
    .A2(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[12][1] ),
    .X(_10672_));
 sky130_fd_sc_hd__a21bo_1 _18203_ (.A1(_10608_),
    .A2(_10645_),
    .B1_N(_10672_),
    .X(_10673_));
 sky130_fd_sc_hd__xor2_2 _18204_ (.A(_10671_),
    .B(_10673_),
    .X(_10674_));
 sky130_fd_sc_hd__xor2_2 _18205_ (.A(_10670_),
    .B(_10674_),
    .X(_10675_));
 sky130_fd_sc_hd__or2_1 _18206_ (.A(_10647_),
    .B(_10654_),
    .X(_10676_));
 sky130_fd_sc_hd__o21ai_2 _18207_ (.A1(_10652_),
    .A2(_10653_),
    .B1(_10676_),
    .Y(_10677_));
 sky130_fd_sc_hd__xor2_2 _18208_ (.A(_10675_),
    .B(_10677_),
    .X(_10678_));
 sky130_fd_sc_hd__nand2_1 _18209_ (.A(_10656_),
    .B(_10659_),
    .Y(_10679_));
 sky130_fd_sc_hd__nor2_1 _18210_ (.A(_10678_),
    .B(_10679_),
    .Y(_10680_));
 sky130_fd_sc_hd__a21o_1 _18211_ (.A1(_10678_),
    .A2(_10679_),
    .B1(_09292_),
    .X(_10681_));
 sky130_fd_sc_hd__o221a_1 _18212_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[4] ),
    .A2(_10364_),
    .B1(_10680_),
    .B2(_10681_),
    .C1(_09886_),
    .X(_00652_));
 sky130_fd_sc_hd__nor2_1 _18213_ (.A(_10659_),
    .B(_10678_),
    .Y(_10682_));
 sky130_fd_sc_hd__and2b_1 _18214_ (.A_N(_10670_),
    .B(_10674_),
    .X(_10683_));
 sky130_fd_sc_hd__nand2_1 _18215_ (.A(_10577_),
    .B(_10610_),
    .Y(_10684_));
 sky130_fd_sc_hd__nand2_1 _18216_ (.A(_10585_),
    .B(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[2] ),
    .Y(_10685_));
 sky130_fd_sc_hd__and3_1 _18217_ (.A(\top_inst.grid_inst.data_path_wires[12][2] ),
    .B(\top_inst.grid_inst.data_path_wires[12][1] ),
    .C(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[4] ),
    .X(_10686_));
 sky130_fd_sc_hd__a22o_1 _18218_ (.A1(\top_inst.grid_inst.data_path_wires[12][1] ),
    .A2(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[12][2] ),
    .X(_10687_));
 sky130_fd_sc_hd__a21bo_1 _18219_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[3] ),
    .A2(_10686_),
    .B1_N(_10687_),
    .X(_10688_));
 sky130_fd_sc_hd__xor2_2 _18220_ (.A(_10685_),
    .B(_10688_),
    .X(_10689_));
 sky130_fd_sc_hd__xnor2_2 _18221_ (.A(_10684_),
    .B(_10689_),
    .Y(_10690_));
 sky130_fd_sc_hd__a21boi_2 _18222_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[4] ),
    .A2(_10664_),
    .B1_N(_10665_),
    .Y(_10691_));
 sky130_fd_sc_hd__a32o_1 _18223_ (.A1(_10581_),
    .A2(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[2] ),
    .A3(_10672_),
    .B1(_10645_),
    .B2(_10608_),
    .X(_10692_));
 sky130_fd_sc_hd__a22o_1 _18224_ (.A1(\top_inst.grid_inst.data_path_wires[12][4] ),
    .A2(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[12][5] ),
    .X(_10693_));
 sky130_fd_sc_hd__nand4_1 _18225_ (.A(\top_inst.grid_inst.data_path_wires[12][5] ),
    .B(\top_inst.grid_inst.data_path_wires[12][4] ),
    .C(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[0] ),
    .Y(_10694_));
 sky130_fd_sc_hd__nand2_1 _18226_ (.A(_10693_),
    .B(_10694_),
    .Y(_10695_));
 sky130_fd_sc_hd__xor2_2 _18227_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[5] ),
    .B(_10695_),
    .X(_10696_));
 sky130_fd_sc_hd__xnor2_2 _18228_ (.A(_10692_),
    .B(_10696_),
    .Y(_10697_));
 sky130_fd_sc_hd__xnor2_2 _18229_ (.A(_10691_),
    .B(_10697_),
    .Y(_10698_));
 sky130_fd_sc_hd__xor2_2 _18230_ (.A(_10690_),
    .B(_10698_),
    .X(_10699_));
 sky130_fd_sc_hd__xor2_2 _18231_ (.A(_10683_),
    .B(_10699_),
    .X(_10700_));
 sky130_fd_sc_hd__nor2_1 _18232_ (.A(_10646_),
    .B(_10667_),
    .Y(_10701_));
 sky130_fd_sc_hd__a21o_1 _18233_ (.A1(_10668_),
    .A2(_10669_),
    .B1(_10701_),
    .X(_10702_));
 sky130_fd_sc_hd__xnor2_2 _18234_ (.A(_10700_),
    .B(_10702_),
    .Y(_10703_));
 sky130_fd_sc_hd__or2b_1 _18235_ (.A(_10675_),
    .B_N(_10677_),
    .X(_10704_));
 sky130_fd_sc_hd__o21a_1 _18236_ (.A1(_10656_),
    .A2(_10678_),
    .B1(_10704_),
    .X(_10705_));
 sky130_fd_sc_hd__xor2_1 _18237_ (.A(_10703_),
    .B(_10705_),
    .X(_10706_));
 sky130_fd_sc_hd__nand2_1 _18238_ (.A(_10682_),
    .B(_10706_),
    .Y(_10707_));
 sky130_fd_sc_hd__o21a_1 _18239_ (.A1(_10682_),
    .A2(_10706_),
    .B1(_08265_),
    .X(_10708_));
 sky130_fd_sc_hd__a22o_1 _18240_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[5] ),
    .A2(_09496_),
    .B1(_10707_),
    .B2(_10708_),
    .X(_10709_));
 sky130_fd_sc_hd__and2_1 _18241_ (.A(_10641_),
    .B(_10709_),
    .X(_10710_));
 sky130_fd_sc_hd__clkbuf_1 _18242_ (.A(_10710_),
    .X(_00653_));
 sky130_fd_sc_hd__nand2_1 _18243_ (.A(_10683_),
    .B(_10699_),
    .Y(_10711_));
 sky130_fd_sc_hd__nand2_1 _18244_ (.A(_10700_),
    .B(_10702_),
    .Y(_10712_));
 sky130_fd_sc_hd__or2b_1 _18245_ (.A(_10696_),
    .B_N(_10692_),
    .X(_10713_));
 sky130_fd_sc_hd__or2b_1 _18246_ (.A(_10691_),
    .B_N(_10697_),
    .X(_10714_));
 sky130_fd_sc_hd__and2_1 _18247_ (.A(_10690_),
    .B(_10698_),
    .X(_10715_));
 sky130_fd_sc_hd__a21boi_1 _18248_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[5] ),
    .A2(_10693_),
    .B1_N(_10694_),
    .Y(_10716_));
 sky130_fd_sc_hd__o2bb2a_1 _18249_ (.A1_N(_10604_),
    .A2_N(_10686_),
    .B1(_10688_),
    .B2(_10685_),
    .X(_10717_));
 sky130_fd_sc_hd__a22o_1 _18250_ (.A1(\top_inst.grid_inst.data_path_wires[12][5] ),
    .A2(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[0] ),
    .B2(_10591_),
    .X(_10718_));
 sky130_fd_sc_hd__nand4_1 _18251_ (.A(_10591_),
    .B(\top_inst.grid_inst.data_path_wires[12][5] ),
    .C(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[0] ),
    .Y(_10719_));
 sky130_fd_sc_hd__nand2_1 _18252_ (.A(_10718_),
    .B(_10719_),
    .Y(_10720_));
 sky130_fd_sc_hd__xor2_1 _18253_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[6] ),
    .B(_10720_),
    .X(_10721_));
 sky130_fd_sc_hd__xor2_1 _18254_ (.A(_10717_),
    .B(_10721_),
    .X(_10722_));
 sky130_fd_sc_hd__xnor2_1 _18255_ (.A(_10716_),
    .B(_10722_),
    .Y(_10723_));
 sky130_fd_sc_hd__or2b_1 _18256_ (.A(_10684_),
    .B_N(_10689_),
    .X(_10724_));
 sky130_fd_sc_hd__a22oi_1 _18257_ (.A1(_10577_),
    .A2(_10612_),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[5] ),
    .B2(_10599_),
    .Y(_10725_));
 sky130_fd_sc_hd__and4_2 _18258_ (.A(_10599_),
    .B(\top_inst.grid_inst.data_path_wires[12][0] ),
    .C(_10612_),
    .D(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[5] ),
    .X(_10726_));
 sky130_fd_sc_hd__nor2_1 _18259_ (.A(_10725_),
    .B(_10726_),
    .Y(_10727_));
 sky130_fd_sc_hd__a22oi_1 _18260_ (.A1(\top_inst.grid_inst.data_path_wires[12][2] ),
    .A2(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[12][3] ),
    .Y(_10728_));
 sky130_fd_sc_hd__and4_1 _18261_ (.A(\top_inst.grid_inst.data_path_wires[12][3] ),
    .B(\top_inst.grid_inst.data_path_wires[12][2] ),
    .C(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[3] ),
    .X(_10729_));
 sky130_fd_sc_hd__and4bb_1 _18262_ (.A_N(_10728_),
    .B_N(_10729_),
    .C(_10606_),
    .D(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[2] ),
    .X(_10730_));
 sky130_fd_sc_hd__o2bb2a_1 _18263_ (.A1_N(_10606_),
    .A2_N(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[2] ),
    .B1(_10728_),
    .B2(_10729_),
    .X(_10731_));
 sky130_fd_sc_hd__nor2_1 _18264_ (.A(_10730_),
    .B(_10731_),
    .Y(_10732_));
 sky130_fd_sc_hd__xnor2_1 _18265_ (.A(_10727_),
    .B(_10732_),
    .Y(_10733_));
 sky130_fd_sc_hd__xor2_1 _18266_ (.A(_10724_),
    .B(_10733_),
    .X(_10734_));
 sky130_fd_sc_hd__nand2_1 _18267_ (.A(_10723_),
    .B(_10734_),
    .Y(_10735_));
 sky130_fd_sc_hd__or2_1 _18268_ (.A(_10723_),
    .B(_10734_),
    .X(_10736_));
 sky130_fd_sc_hd__and3_1 _18269_ (.A(_10715_),
    .B(_10735_),
    .C(_10736_),
    .X(_10737_));
 sky130_fd_sc_hd__a21oi_1 _18270_ (.A1(_10735_),
    .A2(_10736_),
    .B1(_10715_),
    .Y(_10738_));
 sky130_fd_sc_hd__a211oi_2 _18271_ (.A1(_10713_),
    .A2(_10714_),
    .B1(_10737_),
    .C1(_10738_),
    .Y(_10739_));
 sky130_fd_sc_hd__o211a_1 _18272_ (.A1(_10737_),
    .A2(_10738_),
    .B1(_10713_),
    .C1(_10714_),
    .X(_10740_));
 sky130_fd_sc_hd__a211o_1 _18273_ (.A1(_10711_),
    .A2(_10712_),
    .B1(_10739_),
    .C1(_10740_),
    .X(_10741_));
 sky130_fd_sc_hd__o211ai_1 _18274_ (.A1(_10739_),
    .A2(_10740_),
    .B1(_10711_),
    .C1(_10712_),
    .Y(_10742_));
 sky130_fd_sc_hd__and4bb_1 _18275_ (.A_N(_10704_),
    .B_N(_10703_),
    .C(_10741_),
    .D(_10742_),
    .X(_10743_));
 sky130_fd_sc_hd__o2bb2a_1 _18276_ (.A1_N(_10741_),
    .A2_N(_10742_),
    .B1(_10704_),
    .B2(_10703_),
    .X(_10744_));
 sky130_fd_sc_hd__nor2_1 _18277_ (.A(_10743_),
    .B(_10744_),
    .Y(_10745_));
 sky130_fd_sc_hd__o31a_1 _18278_ (.A1(_10656_),
    .A2(_10678_),
    .A3(_10703_),
    .B1(_10707_),
    .X(_10746_));
 sky130_fd_sc_hd__xnor2_1 _18279_ (.A(_10745_),
    .B(_10746_),
    .Y(_10747_));
 sky130_fd_sc_hd__mux2_1 _18280_ (.A0(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[6] ),
    .A1(_10747_),
    .S(_08307_),
    .X(_10748_));
 sky130_fd_sc_hd__and2_1 _18281_ (.A(_10641_),
    .B(_10748_),
    .X(_10749_));
 sky130_fd_sc_hd__clkbuf_1 _18282_ (.A(_10749_),
    .X(_00654_));
 sky130_fd_sc_hd__or2b_1 _18283_ (.A(_10716_),
    .B_N(_10722_),
    .X(_10750_));
 sky130_fd_sc_hd__o21ai_1 _18284_ (.A1(_10717_),
    .A2(_10721_),
    .B1(_10750_),
    .Y(_10751_));
 sky130_fd_sc_hd__o21ai_1 _18285_ (.A1(_10724_),
    .A2(_10733_),
    .B1(_10735_),
    .Y(_10752_));
 sky130_fd_sc_hd__a21bo_1 _18286_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[6] ),
    .A2(_10718_),
    .B1_N(_10719_),
    .X(_10753_));
 sky130_fd_sc_hd__nor2_1 _18287_ (.A(_10729_),
    .B(_10730_),
    .Y(_10754_));
 sky130_fd_sc_hd__a22o_1 _18288_ (.A1(_10591_),
    .A2(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[12][7] ),
    .X(_10755_));
 sky130_fd_sc_hd__nand4_1 _18289_ (.A(\top_inst.grid_inst.data_path_wires[12][7] ),
    .B(_10591_),
    .C(_10600_),
    .D(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[0] ),
    .Y(_10756_));
 sky130_fd_sc_hd__nand2_1 _18290_ (.A(_10755_),
    .B(_10756_),
    .Y(_10757_));
 sky130_fd_sc_hd__xor2_1 _18291_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[7] ),
    .B(_10757_),
    .X(_10758_));
 sky130_fd_sc_hd__xor2_1 _18292_ (.A(_10754_),
    .B(_10758_),
    .X(_10759_));
 sky130_fd_sc_hd__xnor2_1 _18293_ (.A(_10753_),
    .B(_10759_),
    .Y(_10760_));
 sky130_fd_sc_hd__and2_1 _18294_ (.A(_10727_),
    .B(_10732_),
    .X(_10761_));
 sky130_fd_sc_hd__a22o_1 _18295_ (.A1(\top_inst.grid_inst.data_path_wires[12][3] ),
    .A2(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[3] ),
    .B2(_10606_),
    .X(_10762_));
 sky130_fd_sc_hd__nand4_2 _18296_ (.A(_10606_),
    .B(_10585_),
    .C(_10608_),
    .D(_10604_),
    .Y(_10763_));
 sky130_fd_sc_hd__a22o_1 _18297_ (.A1(_10589_),
    .A2(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[2] ),
    .B1(_10762_),
    .B2(_10763_),
    .X(_10764_));
 sky130_fd_sc_hd__nand4_1 _18298_ (.A(_10589_),
    .B(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[2] ),
    .C(_10762_),
    .D(_10763_),
    .Y(_10765_));
 sky130_fd_sc_hd__nand2_1 _18299_ (.A(_10764_),
    .B(_10765_),
    .Y(_10766_));
 sky130_fd_sc_hd__nand2_1 _18300_ (.A(\top_inst.grid_inst.data_path_wires[12][2] ),
    .B(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[5] ),
    .Y(_10767_));
 sky130_fd_sc_hd__nand2_1 _18301_ (.A(\top_inst.grid_inst.data_path_wires[12][1] ),
    .B(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[6] ),
    .Y(_10768_));
 sky130_fd_sc_hd__and2b_1 _18302_ (.A_N(\top_inst.grid_inst.data_path_wires[12][0] ),
    .B(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[7] ),
    .X(_10769_));
 sky130_fd_sc_hd__xnor2_2 _18303_ (.A(_10768_),
    .B(_10769_),
    .Y(_10770_));
 sky130_fd_sc_hd__xnor2_2 _18304_ (.A(_10767_),
    .B(_10770_),
    .Y(_10771_));
 sky130_fd_sc_hd__xnor2_2 _18305_ (.A(_10726_),
    .B(_10771_),
    .Y(_10772_));
 sky130_fd_sc_hd__xor2_2 _18306_ (.A(_10766_),
    .B(_10772_),
    .X(_10773_));
 sky130_fd_sc_hd__xnor2_1 _18307_ (.A(_10761_),
    .B(_10773_),
    .Y(_10774_));
 sky130_fd_sc_hd__xnor2_1 _18308_ (.A(_10760_),
    .B(_10774_),
    .Y(_10775_));
 sky130_fd_sc_hd__xor2_1 _18309_ (.A(_10752_),
    .B(_10775_),
    .X(_10776_));
 sky130_fd_sc_hd__xnor2_1 _18310_ (.A(_10751_),
    .B(_10776_),
    .Y(_10777_));
 sky130_fd_sc_hd__nor2_1 _18311_ (.A(_10737_),
    .B(_10739_),
    .Y(_10778_));
 sky130_fd_sc_hd__xnor2_1 _18312_ (.A(_10777_),
    .B(_10778_),
    .Y(_10779_));
 sky130_fd_sc_hd__xnor2_1 _18313_ (.A(_10614_),
    .B(_10779_),
    .Y(_10780_));
 sky130_fd_sc_hd__xor2_1 _18314_ (.A(_10741_),
    .B(_10780_),
    .X(_10781_));
 sky130_fd_sc_hd__o21bai_2 _18315_ (.A1(_10744_),
    .A2(_10746_),
    .B1_N(_10743_),
    .Y(_10782_));
 sky130_fd_sc_hd__nor2_1 _18316_ (.A(_10781_),
    .B(_10782_),
    .Y(_10783_));
 sky130_fd_sc_hd__a21o_1 _18317_ (.A1(_10781_),
    .A2(_10782_),
    .B1(_05353_),
    .X(_10784_));
 sky130_fd_sc_hd__a2bb2o_1 _18318_ (.A1_N(_10783_),
    .A2_N(_10784_),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[7] ),
    .B2(_07816_),
    .X(_10785_));
 sky130_fd_sc_hd__and2_1 _18319_ (.A(_10641_),
    .B(_10785_),
    .X(_10786_));
 sky130_fd_sc_hd__clkbuf_1 _18320_ (.A(_10786_),
    .X(_00655_));
 sky130_fd_sc_hd__nor2_1 _18321_ (.A(_10754_),
    .B(_10758_),
    .Y(_10787_));
 sky130_fd_sc_hd__a21o_1 _18322_ (.A1(_10753_),
    .A2(_10759_),
    .B1(_10787_),
    .X(_10788_));
 sky130_fd_sc_hd__a21boi_1 _18323_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[7] ),
    .A2(_10755_),
    .B1_N(_10756_),
    .Y(_10789_));
 sky130_fd_sc_hd__nand2_1 _18324_ (.A(_10763_),
    .B(_10765_),
    .Y(_10790_));
 sky130_fd_sc_hd__o21ai_2 _18325_ (.A1(_10600_),
    .A2(_10597_),
    .B1(\top_inst.grid_inst.data_path_wires[12][7] ),
    .Y(_10791_));
 sky130_fd_sc_hd__and3_1 _18326_ (.A(\top_inst.grid_inst.data_path_wires[12][7] ),
    .B(_10600_),
    .C(_10597_),
    .X(_10792_));
 sky130_fd_sc_hd__nor2_4 _18327_ (.A(_10791_),
    .B(_10792_),
    .Y(_10793_));
 sky130_fd_sc_hd__xnor2_1 _18328_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[8] ),
    .B(_10793_),
    .Y(_10794_));
 sky130_fd_sc_hd__xnor2_1 _18329_ (.A(_10790_),
    .B(_10794_),
    .Y(_10795_));
 sky130_fd_sc_hd__xnor2_1 _18330_ (.A(_10789_),
    .B(_10795_),
    .Y(_10796_));
 sky130_fd_sc_hd__a22o_1 _18331_ (.A1(_10606_),
    .A2(_10608_),
    .B1(_10604_),
    .B2(_10589_),
    .X(_10797_));
 sky130_fd_sc_hd__nand4_2 _18332_ (.A(_10589_),
    .B(_10606_),
    .C(_10608_),
    .D(_10604_),
    .Y(_10798_));
 sky130_fd_sc_hd__a22o_1 _18333_ (.A1(_10592_),
    .A2(_10602_),
    .B1(_10797_),
    .B2(_10798_),
    .X(_10799_));
 sky130_fd_sc_hd__nand4_2 _18334_ (.A(_10592_),
    .B(_10602_),
    .C(_10797_),
    .D(_10798_),
    .Y(_10800_));
 sky130_fd_sc_hd__nand2_1 _18335_ (.A(_10799_),
    .B(_10800_),
    .Y(_10801_));
 sky130_fd_sc_hd__nand2_1 _18336_ (.A(_10585_),
    .B(_10610_),
    .Y(_10802_));
 sky130_fd_sc_hd__and4_1 _18337_ (.A(\top_inst.grid_inst.data_path_wires[12][2] ),
    .B(_10579_),
    .C(_10614_),
    .D(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[6] ),
    .X(_10803_));
 sky130_fd_sc_hd__a22o_1 _18338_ (.A1(_10579_),
    .A2(_10614_),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[6] ),
    .B2(\top_inst.grid_inst.data_path_wires[12][2] ),
    .X(_10804_));
 sky130_fd_sc_hd__and2b_1 _18339_ (.A_N(_10803_),
    .B(_10804_),
    .X(_10805_));
 sky130_fd_sc_hd__xnor2_1 _18340_ (.A(_10802_),
    .B(_10805_),
    .Y(_10806_));
 sky130_fd_sc_hd__and3_1 _18341_ (.A(_10599_),
    .B(_10612_),
    .C(_10769_),
    .X(_10807_));
 sky130_fd_sc_hd__a31oi_2 _18342_ (.A1(_10581_),
    .A2(_10610_),
    .A3(_10770_),
    .B1(_10807_),
    .Y(_10808_));
 sky130_fd_sc_hd__xnor2_1 _18343_ (.A(_10806_),
    .B(_10808_),
    .Y(_10809_));
 sky130_fd_sc_hd__xnor2_1 _18344_ (.A(_10801_),
    .B(_10809_),
    .Y(_10810_));
 sky130_fd_sc_hd__nand2_1 _18345_ (.A(_10726_),
    .B(_10771_),
    .Y(_10811_));
 sky130_fd_sc_hd__o21a_1 _18346_ (.A1(_10766_),
    .A2(_10772_),
    .B1(_10811_),
    .X(_10812_));
 sky130_fd_sc_hd__xnor2_1 _18347_ (.A(_10810_),
    .B(_10812_),
    .Y(_10813_));
 sky130_fd_sc_hd__xnor2_1 _18348_ (.A(_10796_),
    .B(_10813_),
    .Y(_10814_));
 sky130_fd_sc_hd__nand2_1 _18349_ (.A(_10761_),
    .B(_10773_),
    .Y(_10815_));
 sky130_fd_sc_hd__o21a_1 _18350_ (.A1(_10760_),
    .A2(_10774_),
    .B1(_10815_),
    .X(_10816_));
 sky130_fd_sc_hd__xor2_1 _18351_ (.A(_10814_),
    .B(_10816_),
    .X(_10817_));
 sky130_fd_sc_hd__xnor2_1 _18352_ (.A(_10788_),
    .B(_10817_),
    .Y(_10818_));
 sky130_fd_sc_hd__or2b_1 _18353_ (.A(_10775_),
    .B_N(_10752_),
    .X(_10819_));
 sky130_fd_sc_hd__or2b_1 _18354_ (.A(_10776_),
    .B_N(_10751_),
    .X(_10820_));
 sky130_fd_sc_hd__and2_1 _18355_ (.A(_10819_),
    .B(_10820_),
    .X(_10821_));
 sky130_fd_sc_hd__xnor2_1 _18356_ (.A(_10818_),
    .B(_10821_),
    .Y(_10822_));
 sky130_fd_sc_hd__and2b_1 _18357_ (.A_N(_10778_),
    .B(_10777_),
    .X(_10823_));
 sky130_fd_sc_hd__a21oi_1 _18358_ (.A1(_10614_),
    .A2(_10779_),
    .B1(_10823_),
    .Y(_10824_));
 sky130_fd_sc_hd__nor2_1 _18359_ (.A(_10822_),
    .B(_10824_),
    .Y(_10825_));
 sky130_fd_sc_hd__and2_1 _18360_ (.A(_10822_),
    .B(_10824_),
    .X(_10826_));
 sky130_fd_sc_hd__nor2_1 _18361_ (.A(_10825_),
    .B(_10826_),
    .Y(_10827_));
 sky130_fd_sc_hd__nor2_1 _18362_ (.A(_10741_),
    .B(_10780_),
    .Y(_10828_));
 sky130_fd_sc_hd__a21o_1 _18363_ (.A1(_10781_),
    .A2(_10782_),
    .B1(_10828_),
    .X(_10829_));
 sky130_fd_sc_hd__nand2_1 _18364_ (.A(_10827_),
    .B(_10829_),
    .Y(_10830_));
 sky130_fd_sc_hd__buf_8 _18365_ (.A(_05310_),
    .X(_10831_));
 sky130_fd_sc_hd__o21a_1 _18366_ (.A1(_10827_),
    .A2(_10829_),
    .B1(_10831_),
    .X(_10832_));
 sky130_fd_sc_hd__a22o_1 _18367_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[8] ),
    .A2(_09496_),
    .B1(_10830_),
    .B2(_10832_),
    .X(_10833_));
 sky130_fd_sc_hd__and2_1 _18368_ (.A(_10641_),
    .B(_10833_),
    .X(_10834_));
 sky130_fd_sc_hd__clkbuf_1 _18369_ (.A(_10834_),
    .X(_00656_));
 sky130_fd_sc_hd__nor2_1 _18370_ (.A(_10818_),
    .B(_10821_),
    .Y(_10835_));
 sky130_fd_sc_hd__a21o_1 _18371_ (.A1(_10827_),
    .A2(_10829_),
    .B1(_10825_),
    .X(_10836_));
 sky130_fd_sc_hd__or2b_1 _18372_ (.A(_10794_),
    .B_N(_10790_),
    .X(_10837_));
 sky130_fd_sc_hd__or2b_1 _18373_ (.A(_10789_),
    .B_N(_10795_),
    .X(_10838_));
 sky130_fd_sc_hd__nand2_1 _18374_ (.A(_10837_),
    .B(_10838_),
    .Y(_10839_));
 sky130_fd_sc_hd__clkbuf_4 _18375_ (.A(_10792_),
    .X(_10840_));
 sky130_fd_sc_hd__a21o_1 _18376_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[8] ),
    .A2(_10793_),
    .B1(_10840_),
    .X(_10841_));
 sky130_fd_sc_hd__xnor2_1 _18377_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[9] ),
    .B(_10793_),
    .Y(_10842_));
 sky130_fd_sc_hd__a21oi_1 _18378_ (.A1(_10798_),
    .A2(_10800_),
    .B1(_10842_),
    .Y(_10843_));
 sky130_fd_sc_hd__and3_1 _18379_ (.A(_10798_),
    .B(_10800_),
    .C(_10842_),
    .X(_10844_));
 sky130_fd_sc_hd__nor2_1 _18380_ (.A(_10843_),
    .B(_10844_),
    .Y(_10845_));
 sky130_fd_sc_hd__xor2_1 _18381_ (.A(_10841_),
    .B(_10845_),
    .X(_10846_));
 sky130_fd_sc_hd__or2b_1 _18382_ (.A(_10808_),
    .B_N(_10806_),
    .X(_10847_));
 sky130_fd_sc_hd__or2b_1 _18383_ (.A(_10801_),
    .B_N(_10809_),
    .X(_10848_));
 sky130_fd_sc_hd__a22o_1 _18384_ (.A1(\top_inst.grid_inst.data_path_wires[12][5] ),
    .A2(_10608_),
    .B1(_10604_),
    .B2(_10591_),
    .X(_10849_));
 sky130_fd_sc_hd__and4_1 _18385_ (.A(\top_inst.grid_inst.data_path_wires[12][6] ),
    .B(\top_inst.grid_inst.data_path_wires[12][5] ),
    .C(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[3] ),
    .X(_10850_));
 sky130_fd_sc_hd__inv_2 _18386_ (.A(_10850_),
    .Y(_10851_));
 sky130_fd_sc_hd__and2_1 _18387_ (.A(_10849_),
    .B(_10851_),
    .X(_10852_));
 sky130_fd_sc_hd__nand2_4 _18388_ (.A(_10595_),
    .B(_10602_),
    .Y(_10853_));
 sky130_fd_sc_hd__xor2_1 _18389_ (.A(_10852_),
    .B(_10853_),
    .X(_10854_));
 sky130_fd_sc_hd__nand2_1 _18390_ (.A(_10606_),
    .B(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[5] ),
    .Y(_10855_));
 sky130_fd_sc_hd__and4b_1 _18391_ (.A_N(\top_inst.grid_inst.data_path_wires[12][2] ),
    .B(_10614_),
    .C(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[6] ),
    .D(\top_inst.grid_inst.data_path_wires[12][3] ),
    .X(_10856_));
 sky130_fd_sc_hd__inv_2 _18392_ (.A(_10614_),
    .Y(_10857_));
 sky130_fd_sc_hd__o2bb2a_1 _18393_ (.A1_N(\top_inst.grid_inst.data_path_wires[12][3] ),
    .A2_N(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[6] ),
    .B1(_10857_),
    .B2(\top_inst.grid_inst.data_path_wires[12][2] ),
    .X(_10858_));
 sky130_fd_sc_hd__nor2_1 _18394_ (.A(_10856_),
    .B(_10858_),
    .Y(_10859_));
 sky130_fd_sc_hd__xnor2_1 _18395_ (.A(_10855_),
    .B(_10859_),
    .Y(_10860_));
 sky130_fd_sc_hd__a31oi_2 _18396_ (.A1(_10585_),
    .A2(_10610_),
    .A3(_10804_),
    .B1(_10803_),
    .Y(_10861_));
 sky130_fd_sc_hd__xnor2_1 _18397_ (.A(_10860_),
    .B(_10861_),
    .Y(_10862_));
 sky130_fd_sc_hd__xor2_1 _18398_ (.A(_10854_),
    .B(_10862_),
    .X(_10863_));
 sky130_fd_sc_hd__a21oi_1 _18399_ (.A1(_10847_),
    .A2(_10848_),
    .B1(_10863_),
    .Y(_10864_));
 sky130_fd_sc_hd__and3_1 _18400_ (.A(_10847_),
    .B(_10848_),
    .C(_10863_),
    .X(_10865_));
 sky130_fd_sc_hd__nor2_1 _18401_ (.A(_10864_),
    .B(_10865_),
    .Y(_10866_));
 sky130_fd_sc_hd__xnor2_1 _18402_ (.A(_10846_),
    .B(_10866_),
    .Y(_10867_));
 sky130_fd_sc_hd__and2b_1 _18403_ (.A_N(_10812_),
    .B(_10810_),
    .X(_10868_));
 sky130_fd_sc_hd__a21oi_1 _18404_ (.A1(_10796_),
    .A2(_10813_),
    .B1(_10868_),
    .Y(_10869_));
 sky130_fd_sc_hd__xnor2_1 _18405_ (.A(_10867_),
    .B(_10869_),
    .Y(_10870_));
 sky130_fd_sc_hd__xor2_1 _18406_ (.A(_10839_),
    .B(_10870_),
    .X(_10871_));
 sky130_fd_sc_hd__nor2_1 _18407_ (.A(_10814_),
    .B(_10816_),
    .Y(_10872_));
 sky130_fd_sc_hd__a21oi_1 _18408_ (.A1(_10788_),
    .A2(_10817_),
    .B1(_10872_),
    .Y(_10873_));
 sky130_fd_sc_hd__nor2_1 _18409_ (.A(_10871_),
    .B(_10873_),
    .Y(_10874_));
 sky130_fd_sc_hd__and2_1 _18410_ (.A(_10871_),
    .B(_10873_),
    .X(_10875_));
 sky130_fd_sc_hd__nor2_1 _18411_ (.A(_10874_),
    .B(_10875_),
    .Y(_10876_));
 sky130_fd_sc_hd__xnor2_1 _18412_ (.A(_10836_),
    .B(_10876_),
    .Y(_10877_));
 sky130_fd_sc_hd__nor2_1 _18413_ (.A(_10835_),
    .B(_10877_),
    .Y(_10878_));
 sky130_fd_sc_hd__a21o_1 _18414_ (.A1(_10835_),
    .A2(_10877_),
    .B1(_09292_),
    .X(_10879_));
 sky130_fd_sc_hd__o221a_1 _18415_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[9] ),
    .A2(_10364_),
    .B1(_10878_),
    .B2(_10879_),
    .C1(_09886_),
    .X(_00657_));
 sky130_fd_sc_hd__a21o_1 _18416_ (.A1(_10827_),
    .A2(_10829_),
    .B1(_10876_),
    .X(_10880_));
 sky130_fd_sc_hd__a22o_1 _18417_ (.A1(_10836_),
    .A2(_10876_),
    .B1(_10880_),
    .B2(_10835_),
    .X(_10881_));
 sky130_fd_sc_hd__or2_1 _18418_ (.A(_10867_),
    .B(_10869_),
    .X(_10882_));
 sky130_fd_sc_hd__or2b_1 _18419_ (.A(_10870_),
    .B_N(_10839_),
    .X(_10883_));
 sky130_fd_sc_hd__a21o_1 _18420_ (.A1(_10841_),
    .A2(_10845_),
    .B1(_10843_),
    .X(_10884_));
 sky130_fd_sc_hd__a21o_1 _18421_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[9] ),
    .A2(_10793_),
    .B1(_10840_),
    .X(_10885_));
 sky130_fd_sc_hd__a31o_1 _18422_ (.A1(_10595_),
    .A2(_10602_),
    .A3(_10849_),
    .B1(_10850_),
    .X(_10886_));
 sky130_fd_sc_hd__xnor2_1 _18423_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[10] ),
    .B(_10793_),
    .Y(_10887_));
 sky130_fd_sc_hd__xnor2_1 _18424_ (.A(_10886_),
    .B(_10887_),
    .Y(_10888_));
 sky130_fd_sc_hd__xnor2_1 _18425_ (.A(_10885_),
    .B(_10888_),
    .Y(_10889_));
 sky130_fd_sc_hd__or2b_1 _18426_ (.A(_10861_),
    .B_N(_10860_),
    .X(_10890_));
 sky130_fd_sc_hd__or2b_1 _18427_ (.A(_10854_),
    .B_N(_10862_),
    .X(_10891_));
 sky130_fd_sc_hd__and3_1 _18428_ (.A(\top_inst.grid_inst.data_path_wires[12][7] ),
    .B(_10608_),
    .C(_10604_),
    .X(_10892_));
 sky130_fd_sc_hd__a22o_1 _18429_ (.A1(_10591_),
    .A2(_10608_),
    .B1(_10604_),
    .B2(\top_inst.grid_inst.data_path_wires[12][7] ),
    .X(_10893_));
 sky130_fd_sc_hd__a21bo_1 _18430_ (.A1(_10592_),
    .A2(_10892_),
    .B1_N(_10893_),
    .X(_10894_));
 sky130_fd_sc_hd__xor2_1 _18431_ (.A(_10853_),
    .B(_10894_),
    .X(_10895_));
 sky130_fd_sc_hd__nand2_1 _18432_ (.A(_10589_),
    .B(_10610_),
    .Y(_10896_));
 sky130_fd_sc_hd__and4b_1 _18433_ (.A_N(\top_inst.grid_inst.data_path_wires[12][3] ),
    .B(_10614_),
    .C(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[6] ),
    .D(\top_inst.grid_inst.data_path_wires[12][4] ),
    .X(_10897_));
 sky130_fd_sc_hd__o2bb2a_1 _18434_ (.A1_N(\top_inst.grid_inst.data_path_wires[12][4] ),
    .A2_N(_10612_),
    .B1(_10857_),
    .B2(\top_inst.grid_inst.data_path_wires[12][3] ),
    .X(_10898_));
 sky130_fd_sc_hd__nor2_1 _18435_ (.A(_10897_),
    .B(_10898_),
    .Y(_10899_));
 sky130_fd_sc_hd__xnor2_1 _18436_ (.A(_10896_),
    .B(_10899_),
    .Y(_10900_));
 sky130_fd_sc_hd__o21ba_1 _18437_ (.A1(_10855_),
    .A2(_10858_),
    .B1_N(_10856_),
    .X(_10901_));
 sky130_fd_sc_hd__xnor2_1 _18438_ (.A(_10900_),
    .B(_10901_),
    .Y(_10902_));
 sky130_fd_sc_hd__xnor2_1 _18439_ (.A(_10895_),
    .B(_10902_),
    .Y(_10903_));
 sky130_fd_sc_hd__a21oi_1 _18440_ (.A1(_10890_),
    .A2(_10891_),
    .B1(_10903_),
    .Y(_10904_));
 sky130_fd_sc_hd__and3_1 _18441_ (.A(_10890_),
    .B(_10891_),
    .C(_10903_),
    .X(_10905_));
 sky130_fd_sc_hd__or2_1 _18442_ (.A(_10904_),
    .B(_10905_),
    .X(_10906_));
 sky130_fd_sc_hd__xnor2_1 _18443_ (.A(_10889_),
    .B(_10906_),
    .Y(_10907_));
 sky130_fd_sc_hd__a21oi_1 _18444_ (.A1(_10846_),
    .A2(_10866_),
    .B1(_10864_),
    .Y(_10908_));
 sky130_fd_sc_hd__xnor2_1 _18445_ (.A(_10907_),
    .B(_10908_),
    .Y(_10909_));
 sky130_fd_sc_hd__xor2_1 _18446_ (.A(_10884_),
    .B(_10909_),
    .X(_10910_));
 sky130_fd_sc_hd__a21o_1 _18447_ (.A1(_10882_),
    .A2(_10883_),
    .B1(_10910_),
    .X(_10911_));
 sky130_fd_sc_hd__nand3_1 _18448_ (.A(_10882_),
    .B(_10883_),
    .C(_10910_),
    .Y(_10912_));
 sky130_fd_sc_hd__and2_1 _18449_ (.A(_10911_),
    .B(_10912_),
    .X(_10913_));
 sky130_fd_sc_hd__nand2_1 _18450_ (.A(_10874_),
    .B(_10913_),
    .Y(_10914_));
 sky130_fd_sc_hd__or2_1 _18451_ (.A(_10874_),
    .B(_10913_),
    .X(_10915_));
 sky130_fd_sc_hd__and2_1 _18452_ (.A(_10914_),
    .B(_10915_),
    .X(_10916_));
 sky130_fd_sc_hd__nand2_1 _18453_ (.A(_10881_),
    .B(_10916_),
    .Y(_10917_));
 sky130_fd_sc_hd__or2_1 _18454_ (.A(_10881_),
    .B(_10916_),
    .X(_10918_));
 sky130_fd_sc_hd__and2_1 _18455_ (.A(_10917_),
    .B(_10918_),
    .X(_10919_));
 sky130_fd_sc_hd__or2_1 _18456_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[10] ),
    .B(_10639_),
    .X(_10920_));
 sky130_fd_sc_hd__o211a_1 _18457_ (.A1(_10071_),
    .A2(_10919_),
    .B1(_10920_),
    .C1(_10620_),
    .X(_00658_));
 sky130_fd_sc_hd__or2b_1 _18458_ (.A(_10887_),
    .B_N(_10886_),
    .X(_10921_));
 sky130_fd_sc_hd__a21bo_1 _18459_ (.A1(_10885_),
    .A2(_10888_),
    .B1_N(_10921_),
    .X(_10922_));
 sky130_fd_sc_hd__clkbuf_4 _18460_ (.A(_10793_),
    .X(_10923_));
 sky130_fd_sc_hd__a21o_1 _18461_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[10] ),
    .A2(_10923_),
    .B1(_10840_),
    .X(_10924_));
 sky130_fd_sc_hd__xnor2_1 _18462_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[11] ),
    .B(_10793_),
    .Y(_10925_));
 sky130_fd_sc_hd__a32o_1 _18463_ (.A1(_10595_),
    .A2(_10602_),
    .A3(_10893_),
    .B1(_10892_),
    .B2(_10592_),
    .X(_10926_));
 sky130_fd_sc_hd__and2b_1 _18464_ (.A_N(_10925_),
    .B(_10926_),
    .X(_10927_));
 sky130_fd_sc_hd__and2b_1 _18465_ (.A_N(_10926_),
    .B(_10925_),
    .X(_10928_));
 sky130_fd_sc_hd__nor2_1 _18466_ (.A(_10927_),
    .B(_10928_),
    .Y(_10929_));
 sky130_fd_sc_hd__xnor2_1 _18467_ (.A(_10924_),
    .B(_10929_),
    .Y(_10930_));
 sky130_fd_sc_hd__o21ai_2 _18468_ (.A1(_10608_),
    .A2(_10604_),
    .B1(_10595_),
    .Y(_10931_));
 sky130_fd_sc_hd__nor2_2 _18469_ (.A(_10892_),
    .B(_10931_),
    .Y(_10932_));
 sky130_fd_sc_hd__xnor2_4 _18470_ (.A(_10853_),
    .B(_10932_),
    .Y(_10933_));
 sky130_fd_sc_hd__and4_1 _18471_ (.A(_10589_),
    .B(_10587_),
    .C(_10614_),
    .D(_10612_),
    .X(_10934_));
 sky130_fd_sc_hd__a22o_1 _18472_ (.A1(_10587_),
    .A2(_10614_),
    .B1(_10612_),
    .B2(\top_inst.grid_inst.data_path_wires[12][5] ),
    .X(_10935_));
 sky130_fd_sc_hd__and4b_1 _18473_ (.A_N(_10934_),
    .B(_10935_),
    .C(_10592_),
    .D(_10610_),
    .X(_10936_));
 sky130_fd_sc_hd__inv_2 _18474_ (.A(_10935_),
    .Y(_10937_));
 sky130_fd_sc_hd__o2bb2a_1 _18475_ (.A1_N(_10592_),
    .A2_N(_10610_),
    .B1(_10934_),
    .B2(_10937_),
    .X(_10938_));
 sky130_fd_sc_hd__nor2_1 _18476_ (.A(_10936_),
    .B(_10938_),
    .Y(_10939_));
 sky130_fd_sc_hd__o21ba_1 _18477_ (.A1(_10896_),
    .A2(_10898_),
    .B1_N(_10897_),
    .X(_10940_));
 sky130_fd_sc_hd__xnor2_1 _18478_ (.A(_10939_),
    .B(_10940_),
    .Y(_10941_));
 sky130_fd_sc_hd__xnor2_1 _18479_ (.A(_10933_),
    .B(_10941_),
    .Y(_10942_));
 sky130_fd_sc_hd__or2b_1 _18480_ (.A(_10901_),
    .B_N(_10900_),
    .X(_10943_));
 sky130_fd_sc_hd__a21bo_1 _18481_ (.A1(_10895_),
    .A2(_10902_),
    .B1_N(_10943_),
    .X(_10944_));
 sky130_fd_sc_hd__xor2_1 _18482_ (.A(_10942_),
    .B(_10944_),
    .X(_10945_));
 sky130_fd_sc_hd__xor2_1 _18483_ (.A(_10930_),
    .B(_10945_),
    .X(_10946_));
 sky130_fd_sc_hd__o21bai_1 _18484_ (.A1(_10889_),
    .A2(_10905_),
    .B1_N(_10904_),
    .Y(_10947_));
 sky130_fd_sc_hd__xnor2_1 _18485_ (.A(_10946_),
    .B(_10947_),
    .Y(_10948_));
 sky130_fd_sc_hd__xor2_1 _18486_ (.A(_10922_),
    .B(_10948_),
    .X(_10949_));
 sky130_fd_sc_hd__or2b_1 _18487_ (.A(_10909_),
    .B_N(_10884_),
    .X(_10950_));
 sky130_fd_sc_hd__o21a_1 _18488_ (.A1(_10907_),
    .A2(_10908_),
    .B1(_10950_),
    .X(_10951_));
 sky130_fd_sc_hd__or2_1 _18489_ (.A(_10949_),
    .B(_10951_),
    .X(_10952_));
 sky130_fd_sc_hd__nand2_1 _18490_ (.A(_10949_),
    .B(_10951_),
    .Y(_10953_));
 sky130_fd_sc_hd__and2_1 _18491_ (.A(_10952_),
    .B(_10953_),
    .X(_10954_));
 sky130_fd_sc_hd__xnor2_1 _18492_ (.A(_10911_),
    .B(_10954_),
    .Y(_10955_));
 sky130_fd_sc_hd__a21oi_1 _18493_ (.A1(_10914_),
    .A2(_10917_),
    .B1(_10955_),
    .Y(_10956_));
 sky130_fd_sc_hd__buf_4 _18494_ (.A(_05633_),
    .X(_10957_));
 sky130_fd_sc_hd__a31o_1 _18495_ (.A1(_10914_),
    .A2(_10917_),
    .A3(_10955_),
    .B1(_10957_),
    .X(_10958_));
 sky130_fd_sc_hd__o221a_1 _18496_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[11] ),
    .A2(_10364_),
    .B1(_10956_),
    .B2(_10958_),
    .C1(_09886_),
    .X(_00659_));
 sky130_fd_sc_hd__nand2_1 _18497_ (.A(_10911_),
    .B(_10914_),
    .Y(_10959_));
 sky130_fd_sc_hd__a32o_1 _18498_ (.A1(_10881_),
    .A2(_10916_),
    .A3(_10955_),
    .B1(_10959_),
    .B2(_10954_),
    .X(_10960_));
 sky130_fd_sc_hd__nand2_1 _18499_ (.A(_10946_),
    .B(_10947_),
    .Y(_10961_));
 sky130_fd_sc_hd__or2b_1 _18500_ (.A(_10948_),
    .B_N(_10922_),
    .X(_10962_));
 sky130_fd_sc_hd__a21o_1 _18501_ (.A1(_10924_),
    .A2(_10929_),
    .B1(_10927_),
    .X(_10963_));
 sky130_fd_sc_hd__inv_2 _18502_ (.A(_10963_),
    .Y(_10964_));
 sky130_fd_sc_hd__and2b_1 _18503_ (.A_N(_10942_),
    .B(_10944_),
    .X(_10965_));
 sky130_fd_sc_hd__o21ba_1 _18504_ (.A1(_10930_),
    .A2(_10945_),
    .B1_N(_10965_),
    .X(_10966_));
 sky130_fd_sc_hd__a21o_1 _18505_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[11] ),
    .A2(_10923_),
    .B1(_10840_),
    .X(_10967_));
 sky130_fd_sc_hd__o21ba_1 _18506_ (.A1(_10853_),
    .A2(_10931_),
    .B1_N(_10892_),
    .X(_10968_));
 sky130_fd_sc_hd__clkbuf_4 _18507_ (.A(_10968_),
    .X(_10969_));
 sky130_fd_sc_hd__xnor2_1 _18508_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[12] ),
    .B(_10793_),
    .Y(_10970_));
 sky130_fd_sc_hd__nor2_1 _18509_ (.A(_10969_),
    .B(_10970_),
    .Y(_10971_));
 sky130_fd_sc_hd__and2_1 _18510_ (.A(_10968_),
    .B(_10970_),
    .X(_10972_));
 sky130_fd_sc_hd__nor2_1 _18511_ (.A(_10971_),
    .B(_10972_),
    .Y(_10973_));
 sky130_fd_sc_hd__xnor2_1 _18512_ (.A(_10967_),
    .B(_10973_),
    .Y(_10974_));
 sky130_fd_sc_hd__nand2_1 _18513_ (.A(_10595_),
    .B(_10610_),
    .Y(_10975_));
 sky130_fd_sc_hd__nor2_1 _18514_ (.A(_10589_),
    .B(_10857_),
    .Y(_10976_));
 sky130_fd_sc_hd__and3_1 _18515_ (.A(_10591_),
    .B(_10612_),
    .C(_10976_),
    .X(_10977_));
 sky130_fd_sc_hd__a21oi_1 _18516_ (.A1(_10592_),
    .A2(_10612_),
    .B1(_10976_),
    .Y(_10978_));
 sky130_fd_sc_hd__nor3_1 _18517_ (.A(_10975_),
    .B(_10977_),
    .C(_10978_),
    .Y(_10979_));
 sky130_fd_sc_hd__o21a_1 _18518_ (.A1(_10977_),
    .A2(_10978_),
    .B1(_10975_),
    .X(_10980_));
 sky130_fd_sc_hd__nor2_1 _18519_ (.A(_10979_),
    .B(_10980_),
    .Y(_10981_));
 sky130_fd_sc_hd__nor2_1 _18520_ (.A(_10934_),
    .B(_10936_),
    .Y(_10982_));
 sky130_fd_sc_hd__xnor2_1 _18521_ (.A(_10981_),
    .B(_10982_),
    .Y(_10983_));
 sky130_fd_sc_hd__nand2_1 _18522_ (.A(_10933_),
    .B(_10983_),
    .Y(_10984_));
 sky130_fd_sc_hd__or2_1 _18523_ (.A(_10933_),
    .B(_10983_),
    .X(_10985_));
 sky130_fd_sc_hd__nand2_1 _18524_ (.A(_10984_),
    .B(_10985_),
    .Y(_10986_));
 sky130_fd_sc_hd__or3_1 _18525_ (.A(_10936_),
    .B(_10938_),
    .C(_10940_),
    .X(_10987_));
 sky130_fd_sc_hd__a21bo_1 _18526_ (.A1(_10933_),
    .A2(_10941_),
    .B1_N(_10987_),
    .X(_10988_));
 sky130_fd_sc_hd__xor2_1 _18527_ (.A(_10986_),
    .B(_10988_),
    .X(_10989_));
 sky130_fd_sc_hd__xor2_1 _18528_ (.A(_10974_),
    .B(_10989_),
    .X(_10990_));
 sky130_fd_sc_hd__or2b_1 _18529_ (.A(_10966_),
    .B_N(_10990_),
    .X(_10991_));
 sky130_fd_sc_hd__or2b_1 _18530_ (.A(_10990_),
    .B_N(_10966_),
    .X(_10992_));
 sky130_fd_sc_hd__nand2_1 _18531_ (.A(_10991_),
    .B(_10992_),
    .Y(_10993_));
 sky130_fd_sc_hd__xnor2_1 _18532_ (.A(_10964_),
    .B(_10993_),
    .Y(_10994_));
 sky130_fd_sc_hd__a21oi_1 _18533_ (.A1(_10961_),
    .A2(_10962_),
    .B1(_10994_),
    .Y(_10995_));
 sky130_fd_sc_hd__and3_1 _18534_ (.A(_10961_),
    .B(_10962_),
    .C(_10994_),
    .X(_10996_));
 sky130_fd_sc_hd__nor2_1 _18535_ (.A(_10995_),
    .B(_10996_),
    .Y(_10997_));
 sky130_fd_sc_hd__xnor2_1 _18536_ (.A(_10952_),
    .B(_10997_),
    .Y(_10998_));
 sky130_fd_sc_hd__nand2_1 _18537_ (.A(_10960_),
    .B(_10998_),
    .Y(_10999_));
 sky130_fd_sc_hd__or2_1 _18538_ (.A(_10960_),
    .B(_10998_),
    .X(_11000_));
 sky130_fd_sc_hd__and2_1 _18539_ (.A(_10999_),
    .B(_11000_),
    .X(_11001_));
 sky130_fd_sc_hd__or2_1 _18540_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[12] ),
    .B(_10639_),
    .X(_11002_));
 sky130_fd_sc_hd__o211a_1 _18541_ (.A1(_10071_),
    .A2(_11001_),
    .B1(_11002_),
    .C1(_10620_),
    .X(_00660_));
 sky130_fd_sc_hd__or3_1 _18542_ (.A(_10952_),
    .B(_10995_),
    .C(_10996_),
    .X(_11003_));
 sky130_fd_sc_hd__a21o_1 _18543_ (.A1(_10961_),
    .A2(_10962_),
    .B1(_10994_),
    .X(_11004_));
 sky130_fd_sc_hd__a21o_1 _18544_ (.A1(_10967_),
    .A2(_10973_),
    .B1(_10971_),
    .X(_11005_));
 sky130_fd_sc_hd__a21o_1 _18545_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[12] ),
    .A2(_10923_),
    .B1(_10840_),
    .X(_11006_));
 sky130_fd_sc_hd__xnor2_1 _18546_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[13] ),
    .B(_10923_),
    .Y(_11007_));
 sky130_fd_sc_hd__nor2_1 _18547_ (.A(_10969_),
    .B(_11007_),
    .Y(_11008_));
 sky130_fd_sc_hd__and2_1 _18548_ (.A(_10969_),
    .B(_11007_),
    .X(_11009_));
 sky130_fd_sc_hd__nor2_1 _18549_ (.A(_11008_),
    .B(_11009_),
    .Y(_11010_));
 sky130_fd_sc_hd__xnor2_2 _18550_ (.A(_11006_),
    .B(_11010_),
    .Y(_11011_));
 sky130_fd_sc_hd__or3_1 _18551_ (.A(_10979_),
    .B(_10980_),
    .C(_10982_),
    .X(_11012_));
 sky130_fd_sc_hd__nand2_1 _18552_ (.A(\top_inst.grid_inst.data_path_wires[12][7] ),
    .B(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[6] ),
    .Y(_11013_));
 sky130_fd_sc_hd__or3_1 _18553_ (.A(_10591_),
    .B(_10857_),
    .C(_11013_),
    .X(_11014_));
 sky130_fd_sc_hd__o21ai_1 _18554_ (.A1(_10591_),
    .A2(_10857_),
    .B1(_11013_),
    .Y(_11015_));
 sky130_fd_sc_hd__and2_1 _18555_ (.A(_11014_),
    .B(_11015_),
    .X(_11016_));
 sky130_fd_sc_hd__xnor2_1 _18556_ (.A(_10975_),
    .B(_11016_),
    .Y(_11017_));
 sky130_fd_sc_hd__o21ai_1 _18557_ (.A1(_10977_),
    .A2(_10979_),
    .B1(_11017_),
    .Y(_11018_));
 sky130_fd_sc_hd__or3_1 _18558_ (.A(_10977_),
    .B(_10979_),
    .C(_11017_),
    .X(_11019_));
 sky130_fd_sc_hd__and2_1 _18559_ (.A(_11018_),
    .B(_11019_),
    .X(_11020_));
 sky130_fd_sc_hd__nand2_1 _18560_ (.A(_10933_),
    .B(_11020_),
    .Y(_11021_));
 sky130_fd_sc_hd__or2_1 _18561_ (.A(_10933_),
    .B(_11020_),
    .X(_11022_));
 sky130_fd_sc_hd__nand2_1 _18562_ (.A(_11021_),
    .B(_11022_),
    .Y(_11023_));
 sky130_fd_sc_hd__a21o_1 _18563_ (.A1(_11012_),
    .A2(_10984_),
    .B1(_11023_),
    .X(_11024_));
 sky130_fd_sc_hd__nand3_1 _18564_ (.A(_11012_),
    .B(_10984_),
    .C(_11023_),
    .Y(_11025_));
 sky130_fd_sc_hd__nand2_1 _18565_ (.A(_11024_),
    .B(_11025_),
    .Y(_11026_));
 sky130_fd_sc_hd__xor2_2 _18566_ (.A(_11011_),
    .B(_11026_),
    .X(_11027_));
 sky130_fd_sc_hd__or2b_1 _18567_ (.A(_10986_),
    .B_N(_10988_),
    .X(_11028_));
 sky130_fd_sc_hd__o21a_1 _18568_ (.A1(_10974_),
    .A2(_10989_),
    .B1(_11028_),
    .X(_11029_));
 sky130_fd_sc_hd__xor2_1 _18569_ (.A(_11027_),
    .B(_11029_),
    .X(_11030_));
 sky130_fd_sc_hd__xor2_1 _18570_ (.A(_11005_),
    .B(_11030_),
    .X(_11031_));
 sky130_fd_sc_hd__o21a_1 _18571_ (.A1(_10964_),
    .A2(_10993_),
    .B1(_10991_),
    .X(_11032_));
 sky130_fd_sc_hd__or2_1 _18572_ (.A(_11031_),
    .B(_11032_),
    .X(_11033_));
 sky130_fd_sc_hd__nand2_1 _18573_ (.A(_11031_),
    .B(_11032_),
    .Y(_11034_));
 sky130_fd_sc_hd__and2_1 _18574_ (.A(_11033_),
    .B(_11034_),
    .X(_11035_));
 sky130_fd_sc_hd__xnor2_1 _18575_ (.A(_11004_),
    .B(_11035_),
    .Y(_11036_));
 sky130_fd_sc_hd__a21oi_1 _18576_ (.A1(_11003_),
    .A2(_10999_),
    .B1(_11036_),
    .Y(_11037_));
 sky130_fd_sc_hd__a31o_1 _18577_ (.A1(_11003_),
    .A2(_10999_),
    .A3(_11036_),
    .B1(_10957_),
    .X(_11038_));
 sky130_fd_sc_hd__o221a_1 _18578_ (.A1(net1085),
    .A2(_10364_),
    .B1(_11037_),
    .B2(_11038_),
    .C1(_09886_),
    .X(_00661_));
 sky130_fd_sc_hd__nand2_1 _18579_ (.A(_11004_),
    .B(_11003_),
    .Y(_11039_));
 sky130_fd_sc_hd__a32o_1 _18580_ (.A1(_10960_),
    .A2(_10998_),
    .A3(_11036_),
    .B1(_11039_),
    .B2(_11035_),
    .X(_11040_));
 sky130_fd_sc_hd__a21o_1 _18581_ (.A1(_11006_),
    .A2(_11010_),
    .B1(_11008_),
    .X(_11041_));
 sky130_fd_sc_hd__inv_2 _18582_ (.A(_11041_),
    .Y(_11042_));
 sky130_fd_sc_hd__o21a_1 _18583_ (.A1(_11011_),
    .A2(_11026_),
    .B1(_11024_),
    .X(_11043_));
 sky130_fd_sc_hd__a21o_1 _18584_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[13] ),
    .A2(_10923_),
    .B1(_10840_),
    .X(_11044_));
 sky130_fd_sc_hd__and2_1 _18585_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[14] ),
    .B(_10923_),
    .X(_11045_));
 sky130_fd_sc_hd__nor2_1 _18586_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[14] ),
    .B(_10923_),
    .Y(_11046_));
 sky130_fd_sc_hd__or2_1 _18587_ (.A(_11045_),
    .B(_11046_),
    .X(_11047_));
 sky130_fd_sc_hd__xor2_1 _18588_ (.A(_10969_),
    .B(_11047_),
    .X(_11048_));
 sky130_fd_sc_hd__nand2_1 _18589_ (.A(_11044_),
    .B(_11048_),
    .Y(_11049_));
 sky130_fd_sc_hd__or2_1 _18590_ (.A(_11044_),
    .B(_11048_),
    .X(_11050_));
 sky130_fd_sc_hd__nand2_1 _18591_ (.A(_11049_),
    .B(_11050_),
    .Y(_11051_));
 sky130_fd_sc_hd__o211a_1 _18592_ (.A1(_10595_),
    .A2(_10857_),
    .B1(_10975_),
    .C1(_11013_),
    .X(_11052_));
 sky130_fd_sc_hd__and2_1 _18593_ (.A(_10595_),
    .B(_10610_),
    .X(_11053_));
 sky130_fd_sc_hd__nand2_1 _18594_ (.A(_11053_),
    .B(_11016_),
    .Y(_11054_));
 sky130_fd_sc_hd__a22oi_2 _18595_ (.A1(_10612_),
    .A2(_11053_),
    .B1(_11014_),
    .B2(_11054_),
    .Y(_11055_));
 sky130_fd_sc_hd__nor2_1 _18596_ (.A(_11052_),
    .B(_11055_),
    .Y(_11056_));
 sky130_fd_sc_hd__xnor2_1 _18597_ (.A(_10933_),
    .B(_11056_),
    .Y(_11057_));
 sky130_fd_sc_hd__a21oi_1 _18598_ (.A1(_11018_),
    .A2(_11021_),
    .B1(_11057_),
    .Y(_11058_));
 sky130_fd_sc_hd__and3_1 _18599_ (.A(_11018_),
    .B(_11021_),
    .C(_11057_),
    .X(_11059_));
 sky130_fd_sc_hd__nor2_1 _18600_ (.A(_11058_),
    .B(_11059_),
    .Y(_11060_));
 sky130_fd_sc_hd__xnor2_1 _18601_ (.A(_11051_),
    .B(_11060_),
    .Y(_11061_));
 sky130_fd_sc_hd__or2b_1 _18602_ (.A(_11043_),
    .B_N(_11061_),
    .X(_11062_));
 sky130_fd_sc_hd__or2b_1 _18603_ (.A(_11061_),
    .B_N(_11043_),
    .X(_11063_));
 sky130_fd_sc_hd__nand2_1 _18604_ (.A(_11062_),
    .B(_11063_),
    .Y(_11064_));
 sky130_fd_sc_hd__xnor2_2 _18605_ (.A(_11042_),
    .B(_11064_),
    .Y(_11065_));
 sky130_fd_sc_hd__inv_2 _18606_ (.A(_11029_),
    .Y(_11066_));
 sky130_fd_sc_hd__and2b_1 _18607_ (.A_N(_11030_),
    .B(_11005_),
    .X(_11067_));
 sky130_fd_sc_hd__a21oi_2 _18608_ (.A1(_11027_),
    .A2(_11066_),
    .B1(_11067_),
    .Y(_11068_));
 sky130_fd_sc_hd__xor2_2 _18609_ (.A(_11065_),
    .B(_11068_),
    .X(_11069_));
 sky130_fd_sc_hd__xnor2_2 _18610_ (.A(_11033_),
    .B(_11069_),
    .Y(_11070_));
 sky130_fd_sc_hd__xor2_1 _18611_ (.A(_11040_),
    .B(_11070_),
    .X(_11071_));
 sky130_fd_sc_hd__or2_1 _18612_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[14] ),
    .B(_10639_),
    .X(_11072_));
 sky130_fd_sc_hd__o211a_1 _18613_ (.A1(_10071_),
    .A2(_11071_),
    .B1(_11072_),
    .C1(_10620_),
    .X(_00662_));
 sky130_fd_sc_hd__or2b_1 _18614_ (.A(_11033_),
    .B_N(_11069_),
    .X(_11073_));
 sky130_fd_sc_hd__a21boi_1 _18615_ (.A1(_11040_),
    .A2(_11070_),
    .B1_N(_11073_),
    .Y(_11074_));
 sky130_fd_sc_hd__or2_1 _18616_ (.A(_11065_),
    .B(_11068_),
    .X(_11075_));
 sky130_fd_sc_hd__o21ai_1 _18617_ (.A1(_10969_),
    .A2(_11047_),
    .B1(_11049_),
    .Y(_11076_));
 sky130_fd_sc_hd__nor2_1 _18618_ (.A(_10933_),
    .B(_11056_),
    .Y(_11077_));
 sky130_fd_sc_hd__xnor2_1 _18619_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[15] ),
    .B(_10923_),
    .Y(_11078_));
 sky130_fd_sc_hd__nor2_1 _18620_ (.A(_10969_),
    .B(_11078_),
    .Y(_11079_));
 sky130_fd_sc_hd__and2_1 _18621_ (.A(_10969_),
    .B(_11078_),
    .X(_11080_));
 sky130_fd_sc_hd__nor2_1 _18622_ (.A(_11079_),
    .B(_11080_),
    .Y(_11081_));
 sky130_fd_sc_hd__o21a_1 _18623_ (.A1(_10840_),
    .A2(_11045_),
    .B1(_11081_),
    .X(_11082_));
 sky130_fd_sc_hd__nor3_1 _18624_ (.A(_10840_),
    .B(_11045_),
    .C(_11081_),
    .Y(_11083_));
 sky130_fd_sc_hd__or2_1 _18625_ (.A(_11082_),
    .B(_11083_),
    .X(_11084_));
 sky130_fd_sc_hd__xor2_1 _18626_ (.A(_11077_),
    .B(_11084_),
    .X(_11085_));
 sky130_fd_sc_hd__a31o_1 _18627_ (.A1(_11049_),
    .A2(_11050_),
    .A3(_11060_),
    .B1(_11058_),
    .X(_11086_));
 sky130_fd_sc_hd__xnor2_1 _18628_ (.A(_11085_),
    .B(_11086_),
    .Y(_11087_));
 sky130_fd_sc_hd__xor2_1 _18629_ (.A(_11076_),
    .B(_11087_),
    .X(_11088_));
 sky130_fd_sc_hd__o21a_1 _18630_ (.A1(_11042_),
    .A2(_11064_),
    .B1(_11062_),
    .X(_11089_));
 sky130_fd_sc_hd__or2_1 _18631_ (.A(_11088_),
    .B(_11089_),
    .X(_11090_));
 sky130_fd_sc_hd__nand2_1 _18632_ (.A(_11088_),
    .B(_11089_),
    .Y(_11091_));
 sky130_fd_sc_hd__and2_1 _18633_ (.A(_11090_),
    .B(_11091_),
    .X(_11092_));
 sky130_fd_sc_hd__xnor2_1 _18634_ (.A(_11075_),
    .B(_11092_),
    .Y(_11093_));
 sky130_fd_sc_hd__nor2_1 _18635_ (.A(_11074_),
    .B(_11093_),
    .Y(_11094_));
 sky130_fd_sc_hd__a2111o_1 _18636_ (.A1(_11074_),
    .A2(_11093_),
    .B1(_11094_),
    .C1(_05309_),
    .D1(_04861_),
    .X(_11095_));
 sky130_fd_sc_hd__o211a_1 _18637_ (.A1(net1067),
    .A2(_10616_),
    .B1(_11095_),
    .C1(_10620_),
    .X(_00663_));
 sky130_fd_sc_hd__nand2_1 _18638_ (.A(_11075_),
    .B(_11073_),
    .Y(_11096_));
 sky130_fd_sc_hd__a32o_1 _18639_ (.A1(_11040_),
    .A2(_11070_),
    .A3(_11093_),
    .B1(_11096_),
    .B2(_11092_),
    .X(_11097_));
 sky130_fd_sc_hd__inv_2 _18640_ (.A(_10933_),
    .Y(_11098_));
 sky130_fd_sc_hd__o2bb2a_1 _18641_ (.A1_N(_11098_),
    .A2_N(_11055_),
    .B1(_11077_),
    .B2(_11084_),
    .X(_11099_));
 sky130_fd_sc_hd__nand2_1 _18642_ (.A(_11098_),
    .B(_11052_),
    .Y(_11100_));
 sky130_fd_sc_hd__a21o_1 _18643_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[15] ),
    .A2(_10923_),
    .B1(_10840_),
    .X(_11101_));
 sky130_fd_sc_hd__xnor2_2 _18644_ (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[16] ),
    .B(_10923_),
    .Y(_11102_));
 sky130_fd_sc_hd__xor2_1 _18645_ (.A(_10969_),
    .B(_11102_),
    .X(_11103_));
 sky130_fd_sc_hd__xnor2_1 _18646_ (.A(_11101_),
    .B(_11103_),
    .Y(_11104_));
 sky130_fd_sc_hd__xor2_1 _18647_ (.A(_11100_),
    .B(_11104_),
    .X(_11105_));
 sky130_fd_sc_hd__xor2_1 _18648_ (.A(_11099_),
    .B(_11105_),
    .X(_11106_));
 sky130_fd_sc_hd__o21ai_1 _18649_ (.A1(_11079_),
    .A2(_11082_),
    .B1(_11106_),
    .Y(_11107_));
 sky130_fd_sc_hd__or3_1 _18650_ (.A(_11079_),
    .B(_11082_),
    .C(_11106_),
    .X(_11108_));
 sky130_fd_sc_hd__nand2_1 _18651_ (.A(_11107_),
    .B(_11108_),
    .Y(_11109_));
 sky130_fd_sc_hd__and2b_1 _18652_ (.A_N(_11087_),
    .B(_11076_),
    .X(_11110_));
 sky130_fd_sc_hd__a21oi_1 _18653_ (.A1(_11085_),
    .A2(_11086_),
    .B1(_11110_),
    .Y(_11111_));
 sky130_fd_sc_hd__xor2_1 _18654_ (.A(_11109_),
    .B(_11111_),
    .X(_11112_));
 sky130_fd_sc_hd__xnor2_1 _18655_ (.A(_11090_),
    .B(_11112_),
    .Y(_11113_));
 sky130_fd_sc_hd__xor2_1 _18656_ (.A(_11097_),
    .B(_11113_),
    .X(_11114_));
 sky130_fd_sc_hd__or2_1 _18657_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[16] ),
    .B(_10639_),
    .X(_11115_));
 sky130_fd_sc_hd__o211a_1 _18658_ (.A1(_10071_),
    .A2(_11114_),
    .B1(_11115_),
    .C1(_10620_),
    .X(_00664_));
 sky130_fd_sc_hd__buf_2 _18659_ (.A(_05313_),
    .X(_11116_));
 sky130_fd_sc_hd__nor2_1 _18660_ (.A(_11109_),
    .B(_11111_),
    .Y(_11117_));
 sky130_fd_sc_hd__o21a_1 _18661_ (.A1(_11099_),
    .A2(_11105_),
    .B1(_11107_),
    .X(_11118_));
 sky130_fd_sc_hd__a21o_1 _18662_ (.A1(_10969_),
    .A2(_11102_),
    .B1(_11101_),
    .X(_11119_));
 sky130_fd_sc_hd__o21a_1 _18663_ (.A1(_10969_),
    .A2(_11102_),
    .B1(_11119_),
    .X(_11120_));
 sky130_fd_sc_hd__nand2_1 _18664_ (.A(_11100_),
    .B(_11104_),
    .Y(_11121_));
 sky130_fd_sc_hd__o21ba_1 _18665_ (.A1(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[16] ),
    .A2(_10840_),
    .B1_N(_10791_),
    .X(_11122_));
 sky130_fd_sc_hd__xnor2_1 _18666_ (.A(_11121_),
    .B(_11122_),
    .Y(_11123_));
 sky130_fd_sc_hd__xnor2_1 _18667_ (.A(_11120_),
    .B(_11123_),
    .Y(_11124_));
 sky130_fd_sc_hd__xnor2_1 _18668_ (.A(_11118_),
    .B(_11124_),
    .Y(_11125_));
 sky130_fd_sc_hd__xnor2_1 _18669_ (.A(_11117_),
    .B(_11125_),
    .Y(_11126_));
 sky130_fd_sc_hd__and2b_1 _18670_ (.A_N(_11090_),
    .B(_11112_),
    .X(_11127_));
 sky130_fd_sc_hd__a211o_1 _18671_ (.A1(_11097_),
    .A2(_11113_),
    .B1(_11126_),
    .C1(_11127_),
    .X(_11128_));
 sky130_fd_sc_hd__a21oi_1 _18672_ (.A1(_05787_),
    .A2(_11128_),
    .B1(_04867_),
    .Y(_11129_));
 sky130_fd_sc_hd__o21a_1 _18673_ (.A1(net922),
    .A2(_11116_),
    .B1(net167),
    .X(_00665_));
 sky130_fd_sc_hd__o21a_1 _18674_ (.A1(net948),
    .A2(_11116_),
    .B1(net167),
    .X(_00666_));
 sky130_fd_sc_hd__o21a_1 _18675_ (.A1(net939),
    .A2(_11116_),
    .B1(net167),
    .X(_00667_));
 sky130_fd_sc_hd__o21a_1 _18676_ (.A1(net947),
    .A2(_11116_),
    .B1(net167),
    .X(_00668_));
 sky130_fd_sc_hd__o21a_1 _18677_ (.A1(net1046),
    .A2(_11116_),
    .B1(net167),
    .X(_00669_));
 sky130_fd_sc_hd__o21a_1 _18678_ (.A1(net1009),
    .A2(_11116_),
    .B1(net167),
    .X(_00670_));
 sky130_fd_sc_hd__o21a_1 _18679_ (.A1(net949),
    .A2(_11116_),
    .B1(net167),
    .X(_00671_));
 sky130_fd_sc_hd__o21a_1 _18680_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[25] ),
    .A2(_11116_),
    .B1(net167),
    .X(_00672_));
 sky130_fd_sc_hd__o21a_1 _18681_ (.A1(net1028),
    .A2(_11116_),
    .B1(net167),
    .X(_00673_));
 sky130_fd_sc_hd__o21a_1 _18682_ (.A1(net706),
    .A2(_11116_),
    .B1(net167),
    .X(_00674_));
 sky130_fd_sc_hd__clkbuf_4 _18683_ (.A(\top_inst.grid_inst.data_path_wires[13][0] ),
    .X(_11130_));
 sky130_fd_sc_hd__or2_1 _18684_ (.A(_11130_),
    .B(_08674_),
    .X(_11131_));
 sky130_fd_sc_hd__o211a_1 _18685_ (.A1(_10577_),
    .A2(_10584_),
    .B1(_11131_),
    .C1(_10620_),
    .X(_00675_));
 sky130_fd_sc_hd__clkbuf_4 _18686_ (.A(\top_inst.grid_inst.data_path_wires[13][1] ),
    .X(_11132_));
 sky130_fd_sc_hd__buf_2 _18687_ (.A(_06619_),
    .X(_11133_));
 sky130_fd_sc_hd__or2_1 _18688_ (.A(_11132_),
    .B(_11133_),
    .X(_11134_));
 sky130_fd_sc_hd__o211a_1 _18689_ (.A1(_10599_),
    .A2(_10584_),
    .B1(_11134_),
    .C1(_10620_),
    .X(_00676_));
 sky130_fd_sc_hd__clkbuf_4 _18690_ (.A(\top_inst.grid_inst.data_path_wires[13][2] ),
    .X(_11135_));
 sky130_fd_sc_hd__or2_1 _18691_ (.A(_11135_),
    .B(_11133_),
    .X(_11136_));
 sky130_fd_sc_hd__buf_2 _18692_ (.A(_10447_),
    .X(_11137_));
 sky130_fd_sc_hd__o211a_1 _18693_ (.A1(_10581_),
    .A2(_10584_),
    .B1(_11136_),
    .C1(_11137_),
    .X(_00677_));
 sky130_fd_sc_hd__clkbuf_4 _18694_ (.A(\top_inst.grid_inst.data_path_wires[13][3] ),
    .X(_11138_));
 sky130_fd_sc_hd__or2_1 _18695_ (.A(_11138_),
    .B(_11133_),
    .X(_11139_));
 sky130_fd_sc_hd__o211a_1 _18696_ (.A1(_10585_),
    .A2(_10584_),
    .B1(_11139_),
    .C1(_11137_),
    .X(_00678_));
 sky130_fd_sc_hd__clkbuf_4 _18697_ (.A(\top_inst.grid_inst.data_path_wires[13][4] ),
    .X(_11140_));
 sky130_fd_sc_hd__or2_1 _18698_ (.A(_11140_),
    .B(_11133_),
    .X(_11141_));
 sky130_fd_sc_hd__o211a_1 _18699_ (.A1(_10606_),
    .A2(_10584_),
    .B1(_11141_),
    .C1(_11137_),
    .X(_00679_));
 sky130_fd_sc_hd__clkbuf_4 _18700_ (.A(_10583_),
    .X(_11142_));
 sky130_fd_sc_hd__clkbuf_4 _18701_ (.A(\top_inst.grid_inst.data_path_wires[13][5] ),
    .X(_11143_));
 sky130_fd_sc_hd__or2_1 _18702_ (.A(_11143_),
    .B(_11133_),
    .X(_11144_));
 sky130_fd_sc_hd__o211a_1 _18703_ (.A1(_10589_),
    .A2(_11142_),
    .B1(_11144_),
    .C1(_11137_),
    .X(_00680_));
 sky130_fd_sc_hd__buf_2 _18704_ (.A(\top_inst.grid_inst.data_path_wires[13][6] ),
    .X(_11145_));
 sky130_fd_sc_hd__or2_1 _18705_ (.A(_11145_),
    .B(_11133_),
    .X(_11146_));
 sky130_fd_sc_hd__o211a_1 _18706_ (.A1(_10592_),
    .A2(_11142_),
    .B1(_11146_),
    .C1(_11137_),
    .X(_00681_));
 sky130_fd_sc_hd__buf_4 _18707_ (.A(\top_inst.grid_inst.data_path_wires[13][7] ),
    .X(_11147_));
 sky130_fd_sc_hd__or2_1 _18708_ (.A(_11147_),
    .B(_11133_),
    .X(_11148_));
 sky130_fd_sc_hd__o211a_1 _18709_ (.A1(_10595_),
    .A2(_11142_),
    .B1(_11148_),
    .C1(_11137_),
    .X(_00682_));
 sky130_fd_sc_hd__clkbuf_4 _18710_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[0] ),
    .X(_11149_));
 sky130_fd_sc_hd__clkbuf_4 _18711_ (.A(_05772_),
    .X(_11150_));
 sky130_fd_sc_hd__or2_1 _18712_ (.A(_11149_),
    .B(_11150_),
    .X(_11151_));
 sky130_fd_sc_hd__o211a_1 _18713_ (.A1(_11130_),
    .A2(_10607_),
    .B1(_11151_),
    .C1(_11137_),
    .X(_00683_));
 sky130_fd_sc_hd__clkbuf_4 _18714_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[1] ),
    .X(_11152_));
 sky130_fd_sc_hd__or2_1 _18715_ (.A(_11152_),
    .B(_11150_),
    .X(_11153_));
 sky130_fd_sc_hd__o211a_1 _18716_ (.A1(_11132_),
    .A2(_10607_),
    .B1(_11153_),
    .C1(_11137_),
    .X(_00684_));
 sky130_fd_sc_hd__buf_4 _18717_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[2] ),
    .X(_11154_));
 sky130_fd_sc_hd__or2_1 _18718_ (.A(_11154_),
    .B(_11150_),
    .X(_11155_));
 sky130_fd_sc_hd__o211a_1 _18719_ (.A1(_11135_),
    .A2(_10607_),
    .B1(_11155_),
    .C1(_11137_),
    .X(_00685_));
 sky130_fd_sc_hd__clkbuf_4 _18720_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[3] ),
    .X(_11156_));
 sky130_fd_sc_hd__or2_1 _18721_ (.A(_11156_),
    .B(_11150_),
    .X(_11157_));
 sky130_fd_sc_hd__o211a_1 _18722_ (.A1(_11138_),
    .A2(_10607_),
    .B1(_11157_),
    .C1(_11137_),
    .X(_00686_));
 sky130_fd_sc_hd__clkbuf_4 _18723_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[4] ),
    .X(_11158_));
 sky130_fd_sc_hd__or2_1 _18724_ (.A(_11158_),
    .B(_11150_),
    .X(_11159_));
 sky130_fd_sc_hd__clkbuf_4 _18725_ (.A(_10447_),
    .X(_11160_));
 sky130_fd_sc_hd__o211a_1 _18726_ (.A1(_11140_),
    .A2(_10607_),
    .B1(_11159_),
    .C1(_11160_),
    .X(_00687_));
 sky130_fd_sc_hd__clkbuf_4 _18727_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[5] ),
    .X(_11161_));
 sky130_fd_sc_hd__or2_1 _18728_ (.A(_11161_),
    .B(_11150_),
    .X(_11162_));
 sky130_fd_sc_hd__o211a_1 _18729_ (.A1(_11143_),
    .A2(_10607_),
    .B1(_11162_),
    .C1(_11160_),
    .X(_00688_));
 sky130_fd_sc_hd__buf_4 _18730_ (.A(_05755_),
    .X(_11163_));
 sky130_fd_sc_hd__buf_2 _18731_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[6] ),
    .X(_11164_));
 sky130_fd_sc_hd__or2_1 _18732_ (.A(_11164_),
    .B(_11150_),
    .X(_11165_));
 sky130_fd_sc_hd__o211a_1 _18733_ (.A1(_11145_),
    .A2(_11163_),
    .B1(_11165_),
    .C1(_11160_),
    .X(_00689_));
 sky130_fd_sc_hd__or2_1 _18734_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[7] ),
    .B(_11150_),
    .X(_11166_));
 sky130_fd_sc_hd__o211a_1 _18735_ (.A1(_11147_),
    .A2(_11163_),
    .B1(_11166_),
    .C1(_11160_),
    .X(_00690_));
 sky130_fd_sc_hd__and3_1 _18736_ (.A(_11149_),
    .B(_11130_),
    .C(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[0] ),
    .X(_11167_));
 sky130_fd_sc_hd__a21oi_1 _18737_ (.A1(_11149_),
    .A2(_11130_),
    .B1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[0] ),
    .Y(_11168_));
 sky130_fd_sc_hd__o21ai_2 _18738_ (.A1(_11167_),
    .A2(_11168_),
    .B1(_08181_),
    .Y(_11169_));
 sky130_fd_sc_hd__o211a_1 _18739_ (.A1(net990),
    .A2(_10616_),
    .B1(_11169_),
    .C1(_11160_),
    .X(_00691_));
 sky130_fd_sc_hd__a22o_1 _18740_ (.A1(_11132_),
    .A2(_11149_),
    .B1(_11130_),
    .B2(_11152_),
    .X(_11170_));
 sky130_fd_sc_hd__nand4_2 _18741_ (.A(_11152_),
    .B(_11132_),
    .C(_11149_),
    .D(_11130_),
    .Y(_11171_));
 sky130_fd_sc_hd__nand3_1 _18742_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[1] ),
    .B(_11170_),
    .C(_11171_),
    .Y(_11172_));
 sky130_fd_sc_hd__a21o_1 _18743_ (.A1(_11170_),
    .A2(_11171_),
    .B1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[1] ),
    .X(_11173_));
 sky130_fd_sc_hd__a21o_1 _18744_ (.A1(_11172_),
    .A2(_11173_),
    .B1(_11167_),
    .X(_11174_));
 sky130_fd_sc_hd__nand3_2 _18745_ (.A(_11167_),
    .B(_11172_),
    .C(_11173_),
    .Y(_11175_));
 sky130_fd_sc_hd__a21o_1 _18746_ (.A1(_11174_),
    .A2(_11175_),
    .B1(_06682_),
    .X(_11176_));
 sky130_fd_sc_hd__o211a_1 _18747_ (.A1(net977),
    .A2(_10616_),
    .B1(_11176_),
    .C1(_11160_),
    .X(_00692_));
 sky130_fd_sc_hd__buf_4 _18748_ (.A(_07057_),
    .X(_11177_));
 sky130_fd_sc_hd__nand2_1 _18749_ (.A(_11154_),
    .B(_11130_),
    .Y(_11178_));
 sky130_fd_sc_hd__a22o_1 _18750_ (.A1(_11152_),
    .A2(_11132_),
    .B1(_11149_),
    .B2(_11135_),
    .X(_11179_));
 sky130_fd_sc_hd__nand4_1 _18751_ (.A(_11135_),
    .B(_11152_),
    .C(_11132_),
    .D(_11149_),
    .Y(_11180_));
 sky130_fd_sc_hd__nand2_1 _18752_ (.A(_11179_),
    .B(_11180_),
    .Y(_11181_));
 sky130_fd_sc_hd__xnor2_1 _18753_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[2] ),
    .B(_11181_),
    .Y(_11182_));
 sky130_fd_sc_hd__nand2_1 _18754_ (.A(_11171_),
    .B(_11172_),
    .Y(_11183_));
 sky130_fd_sc_hd__xnor2_1 _18755_ (.A(_11182_),
    .B(_11183_),
    .Y(_11184_));
 sky130_fd_sc_hd__or2_1 _18756_ (.A(_11178_),
    .B(_11184_),
    .X(_11185_));
 sky130_fd_sc_hd__nand2_1 _18757_ (.A(_11178_),
    .B(_11184_),
    .Y(_11186_));
 sky130_fd_sc_hd__and2_1 _18758_ (.A(_11185_),
    .B(_11186_),
    .X(_11187_));
 sky130_fd_sc_hd__xnor2_1 _18759_ (.A(_11175_),
    .B(_11187_),
    .Y(_11188_));
 sky130_fd_sc_hd__or2_1 _18760_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[2] ),
    .B(_10639_),
    .X(_11189_));
 sky130_fd_sc_hd__o211a_1 _18761_ (.A1(_11177_),
    .A2(_11188_),
    .B1(_11189_),
    .C1(_11160_),
    .X(_00693_));
 sky130_fd_sc_hd__and2b_1 _18762_ (.A_N(_11175_),
    .B(_11187_),
    .X(_11190_));
 sky130_fd_sc_hd__nand2_1 _18763_ (.A(_11182_),
    .B(_11183_),
    .Y(_11191_));
 sky130_fd_sc_hd__a22o_1 _18764_ (.A1(_11154_),
    .A2(_11132_),
    .B1(_11130_),
    .B2(_11156_),
    .X(_11192_));
 sky130_fd_sc_hd__nand4_4 _18765_ (.A(_11156_),
    .B(_11154_),
    .C(_11132_),
    .D(_11130_),
    .Y(_11193_));
 sky130_fd_sc_hd__nand2_2 _18766_ (.A(_11192_),
    .B(_11193_),
    .Y(_11194_));
 sky130_fd_sc_hd__a22o_1 _18767_ (.A1(_11135_),
    .A2(_11152_),
    .B1(_11149_),
    .B2(_11138_),
    .X(_11195_));
 sky130_fd_sc_hd__nand4_2 _18768_ (.A(_11138_),
    .B(_11135_),
    .C(_11152_),
    .D(_11149_),
    .Y(_11196_));
 sky130_fd_sc_hd__and3_1 _18769_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[3] ),
    .B(_11195_),
    .C(_11196_),
    .X(_11197_));
 sky130_fd_sc_hd__a21oi_2 _18770_ (.A1(_11195_),
    .A2(_11196_),
    .B1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[3] ),
    .Y(_11198_));
 sky130_fd_sc_hd__or2_1 _18771_ (.A(_11197_),
    .B(_11198_),
    .X(_11199_));
 sky130_fd_sc_hd__a21boi_4 _18772_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[2] ),
    .A2(_11179_),
    .B1_N(_11180_),
    .Y(_11200_));
 sky130_fd_sc_hd__xnor2_2 _18773_ (.A(_11199_),
    .B(_11200_),
    .Y(_11201_));
 sky130_fd_sc_hd__xnor2_1 _18774_ (.A(_11194_),
    .B(_11201_),
    .Y(_11202_));
 sky130_fd_sc_hd__a21o_1 _18775_ (.A1(_11191_),
    .A2(_11185_),
    .B1(_11202_),
    .X(_11203_));
 sky130_fd_sc_hd__nand3_1 _18776_ (.A(_11191_),
    .B(_11185_),
    .C(_11202_),
    .Y(_11204_));
 sky130_fd_sc_hd__nand3_1 _18777_ (.A(_11190_),
    .B(_11203_),
    .C(_11204_),
    .Y(_11205_));
 sky130_fd_sc_hd__a21o_1 _18778_ (.A1(_11203_),
    .A2(_11204_),
    .B1(_11190_),
    .X(_11206_));
 sky130_fd_sc_hd__and2_1 _18779_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[3] ),
    .B(_05730_),
    .X(_11207_));
 sky130_fd_sc_hd__a31o_1 _18780_ (.A1(_05887_),
    .A2(_11205_),
    .A3(_11206_),
    .B1(_11207_),
    .X(_11208_));
 sky130_fd_sc_hd__and2_1 _18781_ (.A(_10641_),
    .B(_11208_),
    .X(_11209_));
 sky130_fd_sc_hd__clkbuf_1 _18782_ (.A(_11209_),
    .X(_00694_));
 sky130_fd_sc_hd__a22o_1 _18783_ (.A1(\top_inst.grid_inst.data_path_wires[13][3] ),
    .A2(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[13][4] ),
    .X(_11210_));
 sky130_fd_sc_hd__nand4_1 _18784_ (.A(_11140_),
    .B(_11138_),
    .C(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[0] ),
    .Y(_11211_));
 sky130_fd_sc_hd__nand2_2 _18785_ (.A(_11210_),
    .B(_11211_),
    .Y(_11212_));
 sky130_fd_sc_hd__xor2_4 _18786_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[4] ),
    .B(_11212_),
    .X(_11213_));
 sky130_fd_sc_hd__xor2_2 _18787_ (.A(_11193_),
    .B(_11213_),
    .X(_11214_));
 sky130_fd_sc_hd__a21bo_1 _18788_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[3] ),
    .A2(_11195_),
    .B1_N(_11196_),
    .X(_11215_));
 sky130_fd_sc_hd__xnor2_2 _18789_ (.A(_11214_),
    .B(_11215_),
    .Y(_11216_));
 sky130_fd_sc_hd__nand2_2 _18790_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[2] ),
    .B(_11135_),
    .Y(_11217_));
 sky130_fd_sc_hd__nand4_1 _18791_ (.A(_11158_),
    .B(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[3] ),
    .C(\top_inst.grid_inst.data_path_wires[13][1] ),
    .D(\top_inst.grid_inst.data_path_wires[13][0] ),
    .Y(_11218_));
 sky130_fd_sc_hd__a22o_1 _18792_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[3] ),
    .A2(\top_inst.grid_inst.data_path_wires[13][1] ),
    .B1(\top_inst.grid_inst.data_path_wires[13][0] ),
    .B2(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[4] ),
    .X(_11219_));
 sky130_fd_sc_hd__nand2_1 _18793_ (.A(_11218_),
    .B(_11219_),
    .Y(_11220_));
 sky130_fd_sc_hd__xor2_2 _18794_ (.A(_11217_),
    .B(_11220_),
    .X(_11221_));
 sky130_fd_sc_hd__xnor2_2 _18795_ (.A(_11216_),
    .B(_11221_),
    .Y(_11222_));
 sky130_fd_sc_hd__o32ai_4 _18796_ (.A1(_11197_),
    .A2(_11198_),
    .A3(_11200_),
    .B1(_11201_),
    .B2(_11194_),
    .Y(_11223_));
 sky130_fd_sc_hd__xnor2_2 _18797_ (.A(_11222_),
    .B(_11223_),
    .Y(_11224_));
 sky130_fd_sc_hd__nand2_1 _18798_ (.A(_11203_),
    .B(_11205_),
    .Y(_11225_));
 sky130_fd_sc_hd__nor2_1 _18799_ (.A(_11224_),
    .B(_11225_),
    .Y(_11226_));
 sky130_fd_sc_hd__a21o_1 _18800_ (.A1(_11224_),
    .A2(_11225_),
    .B1(_09292_),
    .X(_11227_));
 sky130_fd_sc_hd__buf_4 _18801_ (.A(_07707_),
    .X(_11228_));
 sky130_fd_sc_hd__o221a_1 _18802_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[4] ),
    .A2(_10364_),
    .B1(_11226_),
    .B2(_11227_),
    .C1(_11228_),
    .X(_00695_));
 sky130_fd_sc_hd__nor2_1 _18803_ (.A(_11205_),
    .B(_11224_),
    .Y(_11229_));
 sky130_fd_sc_hd__and2b_1 _18804_ (.A_N(_11216_),
    .B(_11221_),
    .X(_11230_));
 sky130_fd_sc_hd__nand2_1 _18805_ (.A(_11161_),
    .B(_11130_),
    .Y(_11231_));
 sky130_fd_sc_hd__nand2_1 _18806_ (.A(_11138_),
    .B(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[2] ),
    .Y(_11232_));
 sky130_fd_sc_hd__a22o_1 _18807_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[3] ),
    .A2(\top_inst.grid_inst.data_path_wires[13][2] ),
    .B1(\top_inst.grid_inst.data_path_wires[13][1] ),
    .B2(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[4] ),
    .X(_11233_));
 sky130_fd_sc_hd__nand4_1 _18808_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[3] ),
    .C(\top_inst.grid_inst.data_path_wires[13][2] ),
    .D(\top_inst.grid_inst.data_path_wires[13][1] ),
    .Y(_11234_));
 sky130_fd_sc_hd__nand2_1 _18809_ (.A(_11233_),
    .B(_11234_),
    .Y(_11235_));
 sky130_fd_sc_hd__xor2_2 _18810_ (.A(_11232_),
    .B(_11235_),
    .X(_11236_));
 sky130_fd_sc_hd__xnor2_2 _18811_ (.A(_11231_),
    .B(_11236_),
    .Y(_11237_));
 sky130_fd_sc_hd__a21boi_2 _18812_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[4] ),
    .A2(_11210_),
    .B1_N(_11211_),
    .Y(_11238_));
 sky130_fd_sc_hd__o21ai_2 _18813_ (.A1(_11217_),
    .A2(_11220_),
    .B1(_11218_),
    .Y(_11239_));
 sky130_fd_sc_hd__a22o_1 _18814_ (.A1(\top_inst.grid_inst.data_path_wires[13][4] ),
    .A2(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[13][5] ),
    .X(_11240_));
 sky130_fd_sc_hd__nand4_1 _18815_ (.A(\top_inst.grid_inst.data_path_wires[13][5] ),
    .B(\top_inst.grid_inst.data_path_wires[13][4] ),
    .C(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[0] ),
    .Y(_11241_));
 sky130_fd_sc_hd__nand2_1 _18816_ (.A(_11240_),
    .B(_11241_),
    .Y(_11242_));
 sky130_fd_sc_hd__xor2_2 _18817_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[5] ),
    .B(_11242_),
    .X(_11243_));
 sky130_fd_sc_hd__xnor2_2 _18818_ (.A(_11239_),
    .B(_11243_),
    .Y(_11244_));
 sky130_fd_sc_hd__xnor2_2 _18819_ (.A(_11238_),
    .B(_11244_),
    .Y(_11245_));
 sky130_fd_sc_hd__xor2_2 _18820_ (.A(_11237_),
    .B(_11245_),
    .X(_11246_));
 sky130_fd_sc_hd__xor2_2 _18821_ (.A(_11230_),
    .B(_11246_),
    .X(_11247_));
 sky130_fd_sc_hd__nor2_1 _18822_ (.A(_11193_),
    .B(_11213_),
    .Y(_11248_));
 sky130_fd_sc_hd__a21o_1 _18823_ (.A1(_11214_),
    .A2(_11215_),
    .B1(_11248_),
    .X(_11249_));
 sky130_fd_sc_hd__xnor2_2 _18824_ (.A(_11247_),
    .B(_11249_),
    .Y(_11250_));
 sky130_fd_sc_hd__nand2_1 _18825_ (.A(_11222_),
    .B(_11223_),
    .Y(_11251_));
 sky130_fd_sc_hd__o21ai_1 _18826_ (.A1(_11203_),
    .A2(_11224_),
    .B1(_11251_),
    .Y(_11252_));
 sky130_fd_sc_hd__xnor2_1 _18827_ (.A(_11250_),
    .B(_11252_),
    .Y(_11253_));
 sky130_fd_sc_hd__nand2_1 _18828_ (.A(_11229_),
    .B(_11253_),
    .Y(_11254_));
 sky130_fd_sc_hd__o21a_1 _18829_ (.A1(_11229_),
    .A2(_11253_),
    .B1(_10831_),
    .X(_11255_));
 sky130_fd_sc_hd__a22o_1 _18830_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[5] ),
    .A2(_09496_),
    .B1(_11254_),
    .B2(_11255_),
    .X(_11256_));
 sky130_fd_sc_hd__and2_1 _18831_ (.A(_10641_),
    .B(_11256_),
    .X(_11257_));
 sky130_fd_sc_hd__clkbuf_1 _18832_ (.A(_11257_),
    .X(_00696_));
 sky130_fd_sc_hd__nand2_1 _18833_ (.A(_11230_),
    .B(_11246_),
    .Y(_11258_));
 sky130_fd_sc_hd__nand2_1 _18834_ (.A(_11247_),
    .B(_11249_),
    .Y(_11259_));
 sky130_fd_sc_hd__or2b_1 _18835_ (.A(_11243_),
    .B_N(_11239_),
    .X(_11260_));
 sky130_fd_sc_hd__or2b_1 _18836_ (.A(_11238_),
    .B_N(_11244_),
    .X(_11261_));
 sky130_fd_sc_hd__and2_1 _18837_ (.A(_11237_),
    .B(_11245_),
    .X(_11262_));
 sky130_fd_sc_hd__a21boi_2 _18838_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[5] ),
    .A2(_11240_),
    .B1_N(_11241_),
    .Y(_11263_));
 sky130_fd_sc_hd__o21a_1 _18839_ (.A1(_11232_),
    .A2(_11235_),
    .B1(_11234_),
    .X(_11264_));
 sky130_fd_sc_hd__a22o_1 _18840_ (.A1(\top_inst.grid_inst.data_path_wires[13][5] ),
    .A2(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[13][6] ),
    .X(_11265_));
 sky130_fd_sc_hd__nand4_1 _18841_ (.A(\top_inst.grid_inst.data_path_wires[13][6] ),
    .B(\top_inst.grid_inst.data_path_wires[13][5] ),
    .C(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[1] ),
    .D(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[0] ),
    .Y(_11266_));
 sky130_fd_sc_hd__nand2_1 _18842_ (.A(_11265_),
    .B(_11266_),
    .Y(_11267_));
 sky130_fd_sc_hd__xor2_2 _18843_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[6] ),
    .B(_11267_),
    .X(_11268_));
 sky130_fd_sc_hd__xor2_1 _18844_ (.A(_11264_),
    .B(_11268_),
    .X(_11269_));
 sky130_fd_sc_hd__xnor2_1 _18845_ (.A(_11263_),
    .B(_11269_),
    .Y(_11270_));
 sky130_fd_sc_hd__or2b_1 _18846_ (.A(_11231_),
    .B_N(_11236_),
    .X(_11271_));
 sky130_fd_sc_hd__a22oi_1 _18847_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[5] ),
    .A2(_11132_),
    .B1(\top_inst.grid_inst.data_path_wires[13][0] ),
    .B2(_11164_),
    .Y(_11272_));
 sky130_fd_sc_hd__and4_1 _18848_ (.A(_11164_),
    .B(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[5] ),
    .C(\top_inst.grid_inst.data_path_wires[13][1] ),
    .D(\top_inst.grid_inst.data_path_wires[13][0] ),
    .X(_11273_));
 sky130_fd_sc_hd__nor2_1 _18849_ (.A(_11272_),
    .B(_11273_),
    .Y(_11274_));
 sky130_fd_sc_hd__a22oi_1 _18850_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[3] ),
    .A2(\top_inst.grid_inst.data_path_wires[13][3] ),
    .B1(\top_inst.grid_inst.data_path_wires[13][2] ),
    .B2(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[4] ),
    .Y(_11275_));
 sky130_fd_sc_hd__and4_1 _18851_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[3] ),
    .C(\top_inst.grid_inst.data_path_wires[13][3] ),
    .D(\top_inst.grid_inst.data_path_wires[13][2] ),
    .X(_11276_));
 sky130_fd_sc_hd__and4bb_1 _18852_ (.A_N(_11275_),
    .B_N(_11276_),
    .C(_11140_),
    .D(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[2] ),
    .X(_11277_));
 sky130_fd_sc_hd__o2bb2a_1 _18853_ (.A1_N(_11140_),
    .A2_N(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[2] ),
    .B1(_11275_),
    .B2(_11276_),
    .X(_11278_));
 sky130_fd_sc_hd__nor2_1 _18854_ (.A(_11277_),
    .B(_11278_),
    .Y(_11279_));
 sky130_fd_sc_hd__xnor2_1 _18855_ (.A(_11274_),
    .B(_11279_),
    .Y(_11280_));
 sky130_fd_sc_hd__xor2_1 _18856_ (.A(_11271_),
    .B(_11280_),
    .X(_11281_));
 sky130_fd_sc_hd__nand2_1 _18857_ (.A(_11270_),
    .B(_11281_),
    .Y(_11282_));
 sky130_fd_sc_hd__or2_1 _18858_ (.A(_11270_),
    .B(_11281_),
    .X(_11283_));
 sky130_fd_sc_hd__and3_1 _18859_ (.A(_11262_),
    .B(_11282_),
    .C(_11283_),
    .X(_11284_));
 sky130_fd_sc_hd__a21oi_1 _18860_ (.A1(_11282_),
    .A2(_11283_),
    .B1(_11262_),
    .Y(_11285_));
 sky130_fd_sc_hd__a211oi_2 _18861_ (.A1(_11260_),
    .A2(_11261_),
    .B1(_11284_),
    .C1(_11285_),
    .Y(_11286_));
 sky130_fd_sc_hd__o211a_1 _18862_ (.A1(_11284_),
    .A2(_11285_),
    .B1(_11260_),
    .C1(_11261_),
    .X(_11287_));
 sky130_fd_sc_hd__a211o_1 _18863_ (.A1(_11258_),
    .A2(_11259_),
    .B1(_11286_),
    .C1(_11287_),
    .X(_11288_));
 sky130_fd_sc_hd__o211ai_1 _18864_ (.A1(_11286_),
    .A2(_11287_),
    .B1(_11258_),
    .C1(_11259_),
    .Y(_11289_));
 sky130_fd_sc_hd__and4bb_1 _18865_ (.A_N(_11251_),
    .B_N(_11250_),
    .C(_11288_),
    .D(_11289_),
    .X(_11290_));
 sky130_fd_sc_hd__o2bb2a_1 _18866_ (.A1_N(_11288_),
    .A2_N(_11289_),
    .B1(_11251_),
    .B2(_11250_),
    .X(_11291_));
 sky130_fd_sc_hd__nor2_1 _18867_ (.A(_11290_),
    .B(_11291_),
    .Y(_11292_));
 sky130_fd_sc_hd__o31a_1 _18868_ (.A1(_11203_),
    .A2(_11224_),
    .A3(_11250_),
    .B1(_11254_),
    .X(_11293_));
 sky130_fd_sc_hd__xnor2_1 _18869_ (.A(_11292_),
    .B(_11293_),
    .Y(_11294_));
 sky130_fd_sc_hd__mux2_1 _18870_ (.A0(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[6] ),
    .A1(_11294_),
    .S(_08307_),
    .X(_11295_));
 sky130_fd_sc_hd__and2_1 _18871_ (.A(_10641_),
    .B(_11295_),
    .X(_11296_));
 sky130_fd_sc_hd__clkbuf_1 _18872_ (.A(_11296_),
    .X(_00697_));
 sky130_fd_sc_hd__or2b_1 _18873_ (.A(_11263_),
    .B_N(_11269_),
    .X(_11297_));
 sky130_fd_sc_hd__o21ai_2 _18874_ (.A1(_11264_),
    .A2(_11268_),
    .B1(_11297_),
    .Y(_11298_));
 sky130_fd_sc_hd__o21ai_1 _18875_ (.A1(_11271_),
    .A2(_11280_),
    .B1(_11282_),
    .Y(_11299_));
 sky130_fd_sc_hd__a21bo_1 _18876_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[6] ),
    .A2(_11265_),
    .B1_N(_11266_),
    .X(_11300_));
 sky130_fd_sc_hd__nor2_1 _18877_ (.A(_11276_),
    .B(_11277_),
    .Y(_11301_));
 sky130_fd_sc_hd__a22o_1 _18878_ (.A1(\top_inst.grid_inst.data_path_wires[13][6] ),
    .A2(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[1] ),
    .B1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[13][7] ),
    .X(_11302_));
 sky130_fd_sc_hd__nand4_1 _18879_ (.A(\top_inst.grid_inst.data_path_wires[13][7] ),
    .B(\top_inst.grid_inst.data_path_wires[13][6] ),
    .C(_11152_),
    .D(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[0] ),
    .Y(_11303_));
 sky130_fd_sc_hd__nand2_1 _18880_ (.A(_11302_),
    .B(_11303_),
    .Y(_11304_));
 sky130_fd_sc_hd__xor2_2 _18881_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[7] ),
    .B(_11304_),
    .X(_11305_));
 sky130_fd_sc_hd__xor2_1 _18882_ (.A(_11301_),
    .B(_11305_),
    .X(_11306_));
 sky130_fd_sc_hd__xnor2_1 _18883_ (.A(_11300_),
    .B(_11306_),
    .Y(_11307_));
 sky130_fd_sc_hd__and2_1 _18884_ (.A(_11274_),
    .B(_11279_),
    .X(_11308_));
 sky130_fd_sc_hd__a22o_1 _18885_ (.A1(\top_inst.grid_inst.data_path_wires[13][4] ),
    .A2(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[3] ),
    .B1(_11138_),
    .B2(_11158_),
    .X(_11309_));
 sky130_fd_sc_hd__nand4_2 _18886_ (.A(_11158_),
    .B(\top_inst.grid_inst.data_path_wires[13][4] ),
    .C(_11156_),
    .D(_11138_),
    .Y(_11310_));
 sky130_fd_sc_hd__a22o_1 _18887_ (.A1(_11143_),
    .A2(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[2] ),
    .B1(_11309_),
    .B2(_11310_),
    .X(_11311_));
 sky130_fd_sc_hd__nand4_1 _18888_ (.A(_11143_),
    .B(_11154_),
    .C(_11309_),
    .D(_11310_),
    .Y(_11312_));
 sky130_fd_sc_hd__nand2_1 _18889_ (.A(_11311_),
    .B(_11312_),
    .Y(_11313_));
 sky130_fd_sc_hd__nand2_1 _18890_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[5] ),
    .B(_11135_),
    .Y(_11314_));
 sky130_fd_sc_hd__nand2_1 _18891_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[6] ),
    .B(\top_inst.grid_inst.data_path_wires[13][1] ),
    .Y(_11315_));
 sky130_fd_sc_hd__and2b_1 _18892_ (.A_N(\top_inst.grid_inst.data_path_wires[13][0] ),
    .B(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[7] ),
    .X(_11316_));
 sky130_fd_sc_hd__xnor2_2 _18893_ (.A(_11315_),
    .B(_11316_),
    .Y(_11317_));
 sky130_fd_sc_hd__xnor2_1 _18894_ (.A(_11314_),
    .B(_11317_),
    .Y(_11318_));
 sky130_fd_sc_hd__xnor2_1 _18895_ (.A(_11273_),
    .B(_11318_),
    .Y(_11319_));
 sky130_fd_sc_hd__xor2_1 _18896_ (.A(_11313_),
    .B(_11319_),
    .X(_11320_));
 sky130_fd_sc_hd__xnor2_1 _18897_ (.A(_11308_),
    .B(_11320_),
    .Y(_11321_));
 sky130_fd_sc_hd__xnor2_1 _18898_ (.A(_11307_),
    .B(_11321_),
    .Y(_11322_));
 sky130_fd_sc_hd__xor2_1 _18899_ (.A(_11299_),
    .B(_11322_),
    .X(_11323_));
 sky130_fd_sc_hd__xnor2_1 _18900_ (.A(_11298_),
    .B(_11323_),
    .Y(_11324_));
 sky130_fd_sc_hd__nor2_1 _18901_ (.A(_11284_),
    .B(_11286_),
    .Y(_11325_));
 sky130_fd_sc_hd__xnor2_1 _18902_ (.A(_11324_),
    .B(_11325_),
    .Y(_11326_));
 sky130_fd_sc_hd__xnor2_1 _18903_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[7] ),
    .B(_11326_),
    .Y(_11327_));
 sky130_fd_sc_hd__xor2_1 _18904_ (.A(_11288_),
    .B(_11327_),
    .X(_11328_));
 sky130_fd_sc_hd__o21bai_2 _18905_ (.A1(_11291_),
    .A2(_11293_),
    .B1_N(_11290_),
    .Y(_11329_));
 sky130_fd_sc_hd__nor2_1 _18906_ (.A(_11328_),
    .B(_11329_),
    .Y(_11330_));
 sky130_fd_sc_hd__a21o_1 _18907_ (.A1(_11328_),
    .A2(_11329_),
    .B1(_05353_),
    .X(_11331_));
 sky130_fd_sc_hd__a2bb2o_1 _18908_ (.A1_N(_11330_),
    .A2_N(_11331_),
    .B1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[7] ),
    .B2(_07816_),
    .X(_11332_));
 sky130_fd_sc_hd__and2_1 _18909_ (.A(_10641_),
    .B(_11332_),
    .X(_11333_));
 sky130_fd_sc_hd__clkbuf_1 _18910_ (.A(_11333_),
    .X(_00698_));
 sky130_fd_sc_hd__nor2_1 _18911_ (.A(_11301_),
    .B(_11305_),
    .Y(_11334_));
 sky130_fd_sc_hd__a21o_1 _18912_ (.A1(_11300_),
    .A2(_11306_),
    .B1(_11334_),
    .X(_11335_));
 sky130_fd_sc_hd__a21boi_2 _18913_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[7] ),
    .A2(_11302_),
    .B1_N(_11303_),
    .Y(_11336_));
 sky130_fd_sc_hd__nand2_1 _18914_ (.A(_11310_),
    .B(_11312_),
    .Y(_11337_));
 sky130_fd_sc_hd__o21ai_4 _18915_ (.A1(_11152_),
    .A2(_11149_),
    .B1(_11147_),
    .Y(_11338_));
 sky130_fd_sc_hd__and3_1 _18916_ (.A(\top_inst.grid_inst.data_path_wires[13][7] ),
    .B(_11152_),
    .C(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[0] ),
    .X(_11339_));
 sky130_fd_sc_hd__nor2_4 _18917_ (.A(_11338_),
    .B(_11339_),
    .Y(_11340_));
 sky130_fd_sc_hd__xnor2_1 _18918_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[8] ),
    .B(_11340_),
    .Y(_11341_));
 sky130_fd_sc_hd__xnor2_1 _18919_ (.A(_11337_),
    .B(_11341_),
    .Y(_11342_));
 sky130_fd_sc_hd__xnor2_1 _18920_ (.A(_11336_),
    .B(_11342_),
    .Y(_11343_));
 sky130_fd_sc_hd__a22o_1 _18921_ (.A1(_11158_),
    .A2(_11140_),
    .B1(_11156_),
    .B2(_11143_),
    .X(_11344_));
 sky130_fd_sc_hd__nand4_2 _18922_ (.A(_11143_),
    .B(_11158_),
    .C(_11140_),
    .D(_11156_),
    .Y(_11345_));
 sky130_fd_sc_hd__a22o_1 _18923_ (.A1(_11145_),
    .A2(_11154_),
    .B1(_11344_),
    .B2(_11345_),
    .X(_11346_));
 sky130_fd_sc_hd__nand4_1 _18924_ (.A(_11145_),
    .B(_11154_),
    .C(_11344_),
    .D(_11345_),
    .Y(_11347_));
 sky130_fd_sc_hd__nand2_1 _18925_ (.A(_11346_),
    .B(_11347_),
    .Y(_11348_));
 sky130_fd_sc_hd__nand2_1 _18926_ (.A(_11161_),
    .B(_11138_),
    .Y(_11349_));
 sky130_fd_sc_hd__and4b_1 _18927_ (.A_N(\top_inst.grid_inst.data_path_wires[13][1] ),
    .B(\top_inst.grid_inst.data_path_wires[13][2] ),
    .C(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[6] ),
    .D(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[7] ),
    .X(_11350_));
 sky130_fd_sc_hd__inv_2 _18928_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[7] ),
    .Y(_11351_));
 sky130_fd_sc_hd__a2bb2o_1 _18929_ (.A1_N(_11351_),
    .A2_N(\top_inst.grid_inst.data_path_wires[13][1] ),
    .B1(\top_inst.grid_inst.data_path_wires[13][2] ),
    .B2(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[6] ),
    .X(_11352_));
 sky130_fd_sc_hd__and2b_1 _18930_ (.A_N(_11350_),
    .B(_11352_),
    .X(_11353_));
 sky130_fd_sc_hd__xnor2_1 _18931_ (.A(_11349_),
    .B(_11353_),
    .Y(_11354_));
 sky130_fd_sc_hd__and3_1 _18932_ (.A(_11164_),
    .B(_11132_),
    .C(_11316_),
    .X(_11355_));
 sky130_fd_sc_hd__a31oi_2 _18933_ (.A1(_11161_),
    .A2(_11135_),
    .A3(_11317_),
    .B1(_11355_),
    .Y(_11356_));
 sky130_fd_sc_hd__xnor2_1 _18934_ (.A(_11354_),
    .B(_11356_),
    .Y(_11357_));
 sky130_fd_sc_hd__xnor2_1 _18935_ (.A(_11348_),
    .B(_11357_),
    .Y(_11358_));
 sky130_fd_sc_hd__nand2_1 _18936_ (.A(_11273_),
    .B(_11318_),
    .Y(_11359_));
 sky130_fd_sc_hd__o21a_1 _18937_ (.A1(_11313_),
    .A2(_11319_),
    .B1(_11359_),
    .X(_11360_));
 sky130_fd_sc_hd__xnor2_1 _18938_ (.A(_11358_),
    .B(_11360_),
    .Y(_11361_));
 sky130_fd_sc_hd__xnor2_1 _18939_ (.A(_11343_),
    .B(_11361_),
    .Y(_11362_));
 sky130_fd_sc_hd__nand2_1 _18940_ (.A(_11308_),
    .B(_11320_),
    .Y(_11363_));
 sky130_fd_sc_hd__o21a_1 _18941_ (.A1(_11307_),
    .A2(_11321_),
    .B1(_11363_),
    .X(_11364_));
 sky130_fd_sc_hd__xor2_1 _18942_ (.A(_11362_),
    .B(_11364_),
    .X(_11365_));
 sky130_fd_sc_hd__xnor2_1 _18943_ (.A(_11335_),
    .B(_11365_),
    .Y(_11366_));
 sky130_fd_sc_hd__or2b_1 _18944_ (.A(_11322_),
    .B_N(_11299_),
    .X(_11367_));
 sky130_fd_sc_hd__or2b_1 _18945_ (.A(_11323_),
    .B_N(_11298_),
    .X(_11368_));
 sky130_fd_sc_hd__and2_1 _18946_ (.A(_11367_),
    .B(_11368_),
    .X(_11369_));
 sky130_fd_sc_hd__xnor2_1 _18947_ (.A(_11366_),
    .B(_11369_),
    .Y(_11370_));
 sky130_fd_sc_hd__and2b_1 _18948_ (.A_N(_11325_),
    .B(_11324_),
    .X(_11371_));
 sky130_fd_sc_hd__a21oi_1 _18949_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[7] ),
    .A2(_11326_),
    .B1(_11371_),
    .Y(_11372_));
 sky130_fd_sc_hd__nor2_1 _18950_ (.A(_11370_),
    .B(_11372_),
    .Y(_11373_));
 sky130_fd_sc_hd__and2_1 _18951_ (.A(_11370_),
    .B(_11372_),
    .X(_11374_));
 sky130_fd_sc_hd__nor2_1 _18952_ (.A(_11373_),
    .B(_11374_),
    .Y(_11375_));
 sky130_fd_sc_hd__nor2_1 _18953_ (.A(_11288_),
    .B(_11327_),
    .Y(_11376_));
 sky130_fd_sc_hd__a21o_1 _18954_ (.A1(_11328_),
    .A2(_11329_),
    .B1(_11376_),
    .X(_11377_));
 sky130_fd_sc_hd__nand2_1 _18955_ (.A(_11375_),
    .B(_11377_),
    .Y(_11378_));
 sky130_fd_sc_hd__o21a_1 _18956_ (.A1(_11375_),
    .A2(_11377_),
    .B1(_10831_),
    .X(_11379_));
 sky130_fd_sc_hd__a22o_1 _18957_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[8] ),
    .A2(_09496_),
    .B1(_11378_),
    .B2(_11379_),
    .X(_11380_));
 sky130_fd_sc_hd__and2_1 _18958_ (.A(_10641_),
    .B(_11380_),
    .X(_11381_));
 sky130_fd_sc_hd__clkbuf_1 _18959_ (.A(_11381_),
    .X(_00699_));
 sky130_fd_sc_hd__nor2_1 _18960_ (.A(_11366_),
    .B(_11369_),
    .Y(_11382_));
 sky130_fd_sc_hd__a21o_1 _18961_ (.A1(_11375_),
    .A2(_11377_),
    .B1(_11373_),
    .X(_11383_));
 sky130_fd_sc_hd__or2b_1 _18962_ (.A(_11341_),
    .B_N(_11337_),
    .X(_11384_));
 sky130_fd_sc_hd__or2b_1 _18963_ (.A(_11336_),
    .B_N(_11342_),
    .X(_11385_));
 sky130_fd_sc_hd__nand2_1 _18964_ (.A(_11384_),
    .B(_11385_),
    .Y(_11386_));
 sky130_fd_sc_hd__clkbuf_4 _18965_ (.A(_11339_),
    .X(_11387_));
 sky130_fd_sc_hd__a21o_1 _18966_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[8] ),
    .A2(_11340_),
    .B1(_11387_),
    .X(_11388_));
 sky130_fd_sc_hd__xnor2_1 _18967_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[9] ),
    .B(_11340_),
    .Y(_11389_));
 sky130_fd_sc_hd__a21oi_1 _18968_ (.A1(_11345_),
    .A2(_11347_),
    .B1(_11389_),
    .Y(_11390_));
 sky130_fd_sc_hd__and3_1 _18969_ (.A(_11345_),
    .B(_11347_),
    .C(_11389_),
    .X(_11391_));
 sky130_fd_sc_hd__nor2_1 _18970_ (.A(_11390_),
    .B(_11391_),
    .Y(_11392_));
 sky130_fd_sc_hd__xor2_1 _18971_ (.A(_11388_),
    .B(_11392_),
    .X(_11393_));
 sky130_fd_sc_hd__or2b_1 _18972_ (.A(_11356_),
    .B_N(_11354_),
    .X(_11394_));
 sky130_fd_sc_hd__or2b_1 _18973_ (.A(_11348_),
    .B_N(_11357_),
    .X(_11395_));
 sky130_fd_sc_hd__a22o_1 _18974_ (.A1(\top_inst.grid_inst.data_path_wires[13][5] ),
    .A2(_11158_),
    .B1(_11156_),
    .B2(\top_inst.grid_inst.data_path_wires[13][6] ),
    .X(_11396_));
 sky130_fd_sc_hd__and4_1 _18975_ (.A(\top_inst.grid_inst.data_path_wires[13][6] ),
    .B(\top_inst.grid_inst.data_path_wires[13][5] ),
    .C(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[3] ),
    .X(_11397_));
 sky130_fd_sc_hd__inv_2 _18976_ (.A(_11397_),
    .Y(_11398_));
 sky130_fd_sc_hd__and2_1 _18977_ (.A(_11396_),
    .B(_11398_),
    .X(_11399_));
 sky130_fd_sc_hd__nand2_4 _18978_ (.A(_11147_),
    .B(_11154_),
    .Y(_11400_));
 sky130_fd_sc_hd__xor2_1 _18979_ (.A(_11399_),
    .B(_11400_),
    .X(_11401_));
 sky130_fd_sc_hd__nand2_1 _18980_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[5] ),
    .B(_11140_),
    .Y(_11402_));
 sky130_fd_sc_hd__and4b_1 _18981_ (.A_N(\top_inst.grid_inst.data_path_wires[13][2] ),
    .B(\top_inst.grid_inst.data_path_wires[13][3] ),
    .C(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[6] ),
    .D(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[7] ),
    .X(_11403_));
 sky130_fd_sc_hd__o2bb2a_1 _18982_ (.A1_N(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[6] ),
    .A2_N(\top_inst.grid_inst.data_path_wires[13][3] ),
    .B1(_11135_),
    .B2(_11351_),
    .X(_11404_));
 sky130_fd_sc_hd__nor2_1 _18983_ (.A(_11403_),
    .B(_11404_),
    .Y(_11405_));
 sky130_fd_sc_hd__xnor2_1 _18984_ (.A(_11402_),
    .B(_11405_),
    .Y(_11406_));
 sky130_fd_sc_hd__a31oi_2 _18985_ (.A1(_11161_),
    .A2(_11138_),
    .A3(_11352_),
    .B1(_11350_),
    .Y(_11407_));
 sky130_fd_sc_hd__xnor2_1 _18986_ (.A(_11406_),
    .B(_11407_),
    .Y(_11408_));
 sky130_fd_sc_hd__xor2_1 _18987_ (.A(_11401_),
    .B(_11408_),
    .X(_11409_));
 sky130_fd_sc_hd__a21oi_1 _18988_ (.A1(_11394_),
    .A2(_11395_),
    .B1(_11409_),
    .Y(_11410_));
 sky130_fd_sc_hd__and3_1 _18989_ (.A(_11394_),
    .B(_11395_),
    .C(_11409_),
    .X(_11411_));
 sky130_fd_sc_hd__nor2_1 _18990_ (.A(_11410_),
    .B(_11411_),
    .Y(_11412_));
 sky130_fd_sc_hd__xnor2_1 _18991_ (.A(_11393_),
    .B(_11412_),
    .Y(_11413_));
 sky130_fd_sc_hd__and2b_1 _18992_ (.A_N(_11360_),
    .B(_11358_),
    .X(_11414_));
 sky130_fd_sc_hd__a21oi_1 _18993_ (.A1(_11343_),
    .A2(_11361_),
    .B1(_11414_),
    .Y(_11415_));
 sky130_fd_sc_hd__xnor2_1 _18994_ (.A(_11413_),
    .B(_11415_),
    .Y(_11416_));
 sky130_fd_sc_hd__xor2_1 _18995_ (.A(_11386_),
    .B(_11416_),
    .X(_11417_));
 sky130_fd_sc_hd__nor2_1 _18996_ (.A(_11362_),
    .B(_11364_),
    .Y(_11418_));
 sky130_fd_sc_hd__a21oi_1 _18997_ (.A1(_11335_),
    .A2(_11365_),
    .B1(_11418_),
    .Y(_11419_));
 sky130_fd_sc_hd__nor2_1 _18998_ (.A(_11417_),
    .B(_11419_),
    .Y(_11420_));
 sky130_fd_sc_hd__and2_1 _18999_ (.A(_11417_),
    .B(_11419_),
    .X(_11421_));
 sky130_fd_sc_hd__nor2_1 _19000_ (.A(_11420_),
    .B(_11421_),
    .Y(_11422_));
 sky130_fd_sc_hd__xnor2_1 _19001_ (.A(_11383_),
    .B(_11422_),
    .Y(_11423_));
 sky130_fd_sc_hd__nor2_1 _19002_ (.A(_11382_),
    .B(_11423_),
    .Y(_11424_));
 sky130_fd_sc_hd__a21o_1 _19003_ (.A1(_11382_),
    .A2(_11423_),
    .B1(_09292_),
    .X(_11425_));
 sky130_fd_sc_hd__o221a_1 _19004_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[9] ),
    .A2(_10364_),
    .B1(_11424_),
    .B2(_11425_),
    .C1(_11228_),
    .X(_00700_));
 sky130_fd_sc_hd__a21o_1 _19005_ (.A1(_11375_),
    .A2(_11377_),
    .B1(_11422_),
    .X(_11426_));
 sky130_fd_sc_hd__a22o_1 _19006_ (.A1(_11383_),
    .A2(_11422_),
    .B1(_11426_),
    .B2(_11382_),
    .X(_11427_));
 sky130_fd_sc_hd__or2_1 _19007_ (.A(_11413_),
    .B(_11415_),
    .X(_11428_));
 sky130_fd_sc_hd__or2b_1 _19008_ (.A(_11416_),
    .B_N(_11386_),
    .X(_11429_));
 sky130_fd_sc_hd__a21o_1 _19009_ (.A1(_11388_),
    .A2(_11392_),
    .B1(_11390_),
    .X(_11430_));
 sky130_fd_sc_hd__a21o_1 _19010_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[9] ),
    .A2(_11340_),
    .B1(_11387_),
    .X(_11431_));
 sky130_fd_sc_hd__a31o_1 _19011_ (.A1(_11147_),
    .A2(_11154_),
    .A3(_11396_),
    .B1(_11397_),
    .X(_11432_));
 sky130_fd_sc_hd__xnor2_1 _19012_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[10] ),
    .B(_11340_),
    .Y(_11433_));
 sky130_fd_sc_hd__xnor2_1 _19013_ (.A(_11432_),
    .B(_11433_),
    .Y(_11434_));
 sky130_fd_sc_hd__xnor2_1 _19014_ (.A(_11431_),
    .B(_11434_),
    .Y(_11435_));
 sky130_fd_sc_hd__or2b_1 _19015_ (.A(_11407_),
    .B_N(_11406_),
    .X(_11436_));
 sky130_fd_sc_hd__or2b_1 _19016_ (.A(_11401_),
    .B_N(_11408_),
    .X(_11437_));
 sky130_fd_sc_hd__and3_1 _19017_ (.A(\top_inst.grid_inst.data_path_wires[13][7] ),
    .B(_11158_),
    .C(_11156_),
    .X(_11438_));
 sky130_fd_sc_hd__a22o_1 _19018_ (.A1(\top_inst.grid_inst.data_path_wires[13][6] ),
    .A2(_11158_),
    .B1(_11156_),
    .B2(\top_inst.grid_inst.data_path_wires[13][7] ),
    .X(_11439_));
 sky130_fd_sc_hd__a21bo_1 _19019_ (.A1(_11145_),
    .A2(_11438_),
    .B1_N(_11439_),
    .X(_11440_));
 sky130_fd_sc_hd__xor2_1 _19020_ (.A(_11400_),
    .B(_11440_),
    .X(_11441_));
 sky130_fd_sc_hd__nand2_1 _19021_ (.A(_11161_),
    .B(_11143_),
    .Y(_11442_));
 sky130_fd_sc_hd__and4b_1 _19022_ (.A_N(\top_inst.grid_inst.data_path_wires[13][3] ),
    .B(\top_inst.grid_inst.data_path_wires[13][4] ),
    .C(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[6] ),
    .D(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[7] ),
    .X(_11443_));
 sky130_fd_sc_hd__o2bb2a_1 _19023_ (.A1_N(_11164_),
    .A2_N(\top_inst.grid_inst.data_path_wires[13][4] ),
    .B1(\top_inst.grid_inst.data_path_wires[13][3] ),
    .B2(_11351_),
    .X(_11444_));
 sky130_fd_sc_hd__nor2_1 _19024_ (.A(_11443_),
    .B(_11444_),
    .Y(_11445_));
 sky130_fd_sc_hd__xnor2_1 _19025_ (.A(_11442_),
    .B(_11445_),
    .Y(_11446_));
 sky130_fd_sc_hd__o21ba_1 _19026_ (.A1(_11402_),
    .A2(_11404_),
    .B1_N(_11403_),
    .X(_11447_));
 sky130_fd_sc_hd__xnor2_1 _19027_ (.A(_11446_),
    .B(_11447_),
    .Y(_11448_));
 sky130_fd_sc_hd__xnor2_1 _19028_ (.A(_11441_),
    .B(_11448_),
    .Y(_11449_));
 sky130_fd_sc_hd__a21oi_1 _19029_ (.A1(_11436_),
    .A2(_11437_),
    .B1(_11449_),
    .Y(_11450_));
 sky130_fd_sc_hd__and3_1 _19030_ (.A(_11436_),
    .B(_11437_),
    .C(_11449_),
    .X(_11451_));
 sky130_fd_sc_hd__or2_1 _19031_ (.A(_11450_),
    .B(_11451_),
    .X(_11452_));
 sky130_fd_sc_hd__xnor2_1 _19032_ (.A(_11435_),
    .B(_11452_),
    .Y(_11453_));
 sky130_fd_sc_hd__a21oi_1 _19033_ (.A1(_11393_),
    .A2(_11412_),
    .B1(_11410_),
    .Y(_11454_));
 sky130_fd_sc_hd__xnor2_1 _19034_ (.A(_11453_),
    .B(_11454_),
    .Y(_11455_));
 sky130_fd_sc_hd__xor2_1 _19035_ (.A(_11430_),
    .B(_11455_),
    .X(_11456_));
 sky130_fd_sc_hd__a21o_1 _19036_ (.A1(_11428_),
    .A2(_11429_),
    .B1(_11456_),
    .X(_11457_));
 sky130_fd_sc_hd__nand3_1 _19037_ (.A(_11428_),
    .B(_11429_),
    .C(_11456_),
    .Y(_11458_));
 sky130_fd_sc_hd__and2_1 _19038_ (.A(_11457_),
    .B(_11458_),
    .X(_11459_));
 sky130_fd_sc_hd__nand2_1 _19039_ (.A(_11420_),
    .B(_11459_),
    .Y(_11460_));
 sky130_fd_sc_hd__or2_1 _19040_ (.A(_11420_),
    .B(_11459_),
    .X(_11461_));
 sky130_fd_sc_hd__and2_1 _19041_ (.A(_11460_),
    .B(_11461_),
    .X(_11462_));
 sky130_fd_sc_hd__nand2_1 _19042_ (.A(_11427_),
    .B(_11462_),
    .Y(_11463_));
 sky130_fd_sc_hd__or2_1 _19043_ (.A(_11427_),
    .B(_11462_),
    .X(_11464_));
 sky130_fd_sc_hd__and2_1 _19044_ (.A(_11463_),
    .B(_11464_),
    .X(_11465_));
 sky130_fd_sc_hd__or2_1 _19045_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[10] ),
    .B(_10639_),
    .X(_11466_));
 sky130_fd_sc_hd__o211a_1 _19046_ (.A1(_11177_),
    .A2(_11465_),
    .B1(_11466_),
    .C1(_11160_),
    .X(_00701_));
 sky130_fd_sc_hd__or2b_1 _19047_ (.A(_11433_),
    .B_N(_11432_),
    .X(_11467_));
 sky130_fd_sc_hd__a21bo_1 _19048_ (.A1(_11431_),
    .A2(_11434_),
    .B1_N(_11467_),
    .X(_11468_));
 sky130_fd_sc_hd__clkbuf_4 _19049_ (.A(_11340_),
    .X(_11469_));
 sky130_fd_sc_hd__a21o_1 _19050_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[10] ),
    .A2(_11469_),
    .B1(_11387_),
    .X(_11470_));
 sky130_fd_sc_hd__xnor2_1 _19051_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[11] ),
    .B(_11340_),
    .Y(_11471_));
 sky130_fd_sc_hd__a32o_1 _19052_ (.A1(_11147_),
    .A2(_11154_),
    .A3(_11439_),
    .B1(_11438_),
    .B2(_11145_),
    .X(_11472_));
 sky130_fd_sc_hd__and2b_1 _19053_ (.A_N(_11471_),
    .B(_11472_),
    .X(_11473_));
 sky130_fd_sc_hd__and2b_1 _19054_ (.A_N(_11472_),
    .B(_11471_),
    .X(_11474_));
 sky130_fd_sc_hd__nor2_1 _19055_ (.A(_11473_),
    .B(_11474_),
    .Y(_11475_));
 sky130_fd_sc_hd__xnor2_1 _19056_ (.A(_11470_),
    .B(_11475_),
    .Y(_11476_));
 sky130_fd_sc_hd__o21ai_2 _19057_ (.A1(_11158_),
    .A2(_11156_),
    .B1(_11147_),
    .Y(_11477_));
 sky130_fd_sc_hd__nor2_2 _19058_ (.A(_11438_),
    .B(_11477_),
    .Y(_11478_));
 sky130_fd_sc_hd__xnor2_4 _19059_ (.A(_11400_),
    .B(_11478_),
    .Y(_11479_));
 sky130_fd_sc_hd__and4b_1 _19060_ (.A_N(_11140_),
    .B(_11143_),
    .C(_11164_),
    .D(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[7] ),
    .X(_11480_));
 sky130_fd_sc_hd__a2bb2o_1 _19061_ (.A1_N(_11351_),
    .A2_N(_11140_),
    .B1(_11143_),
    .B2(_11164_),
    .X(_11481_));
 sky130_fd_sc_hd__and4b_1 _19062_ (.A_N(_11480_),
    .B(_11481_),
    .C(_11145_),
    .D(_11161_),
    .X(_11482_));
 sky130_fd_sc_hd__inv_2 _19063_ (.A(_11481_),
    .Y(_11483_));
 sky130_fd_sc_hd__o2bb2a_1 _19064_ (.A1_N(_11145_),
    .A2_N(_11161_),
    .B1(_11480_),
    .B2(_11483_),
    .X(_11484_));
 sky130_fd_sc_hd__nor2_1 _19065_ (.A(_11482_),
    .B(_11484_),
    .Y(_11485_));
 sky130_fd_sc_hd__o21ba_1 _19066_ (.A1(_11442_),
    .A2(_11444_),
    .B1_N(_11443_),
    .X(_11486_));
 sky130_fd_sc_hd__xnor2_1 _19067_ (.A(_11485_),
    .B(_11486_),
    .Y(_11487_));
 sky130_fd_sc_hd__xnor2_1 _19068_ (.A(_11479_),
    .B(_11487_),
    .Y(_11488_));
 sky130_fd_sc_hd__or2b_1 _19069_ (.A(_11447_),
    .B_N(_11446_),
    .X(_11489_));
 sky130_fd_sc_hd__a21bo_1 _19070_ (.A1(_11441_),
    .A2(_11448_),
    .B1_N(_11489_),
    .X(_11490_));
 sky130_fd_sc_hd__xor2_1 _19071_ (.A(_11488_),
    .B(_11490_),
    .X(_11491_));
 sky130_fd_sc_hd__xor2_1 _19072_ (.A(_11476_),
    .B(_11491_),
    .X(_11492_));
 sky130_fd_sc_hd__o21bai_2 _19073_ (.A1(_11435_),
    .A2(_11451_),
    .B1_N(_11450_),
    .Y(_11493_));
 sky130_fd_sc_hd__xnor2_1 _19074_ (.A(_11492_),
    .B(_11493_),
    .Y(_11494_));
 sky130_fd_sc_hd__xor2_1 _19075_ (.A(_11468_),
    .B(_11494_),
    .X(_11495_));
 sky130_fd_sc_hd__or2b_1 _19076_ (.A(_11455_),
    .B_N(_11430_),
    .X(_11496_));
 sky130_fd_sc_hd__o21a_1 _19077_ (.A1(_11453_),
    .A2(_11454_),
    .B1(_11496_),
    .X(_11497_));
 sky130_fd_sc_hd__or2_1 _19078_ (.A(_11495_),
    .B(_11497_),
    .X(_11498_));
 sky130_fd_sc_hd__nand2_1 _19079_ (.A(_11495_),
    .B(_11497_),
    .Y(_11499_));
 sky130_fd_sc_hd__and2_1 _19080_ (.A(_11498_),
    .B(_11499_),
    .X(_11500_));
 sky130_fd_sc_hd__xnor2_1 _19081_ (.A(_11457_),
    .B(_11500_),
    .Y(_11501_));
 sky130_fd_sc_hd__a21oi_1 _19082_ (.A1(_11460_),
    .A2(_11463_),
    .B1(_11501_),
    .Y(_11502_));
 sky130_fd_sc_hd__a31o_1 _19083_ (.A1(_11460_),
    .A2(_11463_),
    .A3(_11501_),
    .B1(_10957_),
    .X(_11503_));
 sky130_fd_sc_hd__o221a_1 _19084_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[11] ),
    .A2(_10364_),
    .B1(_11502_),
    .B2(_11503_),
    .C1(_11228_),
    .X(_00702_));
 sky130_fd_sc_hd__nand2_1 _19085_ (.A(_11457_),
    .B(_11460_),
    .Y(_11504_));
 sky130_fd_sc_hd__a32o_1 _19086_ (.A1(_11427_),
    .A2(_11462_),
    .A3(_11501_),
    .B1(_11504_),
    .B2(_11500_),
    .X(_11505_));
 sky130_fd_sc_hd__nand2_1 _19087_ (.A(_11492_),
    .B(_11493_),
    .Y(_11506_));
 sky130_fd_sc_hd__or2b_1 _19088_ (.A(_11494_),
    .B_N(_11468_),
    .X(_11507_));
 sky130_fd_sc_hd__a21o_1 _19089_ (.A1(_11470_),
    .A2(_11475_),
    .B1(_11473_),
    .X(_11508_));
 sky130_fd_sc_hd__inv_2 _19090_ (.A(_11508_),
    .Y(_11509_));
 sky130_fd_sc_hd__and2b_1 _19091_ (.A_N(_11488_),
    .B(_11490_),
    .X(_11510_));
 sky130_fd_sc_hd__o21ba_1 _19092_ (.A1(_11476_),
    .A2(_11491_),
    .B1_N(_11510_),
    .X(_11511_));
 sky130_fd_sc_hd__a21o_1 _19093_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[11] ),
    .A2(_11469_),
    .B1(_11387_),
    .X(_11512_));
 sky130_fd_sc_hd__o21ba_1 _19094_ (.A1(_11400_),
    .A2(_11477_),
    .B1_N(_11438_),
    .X(_11513_));
 sky130_fd_sc_hd__clkbuf_4 _19095_ (.A(_11513_),
    .X(_11514_));
 sky130_fd_sc_hd__xnor2_1 _19096_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[12] ),
    .B(_11340_),
    .Y(_11515_));
 sky130_fd_sc_hd__nor2_1 _19097_ (.A(_11514_),
    .B(_11515_),
    .Y(_11516_));
 sky130_fd_sc_hd__and2_1 _19098_ (.A(_11513_),
    .B(_11515_),
    .X(_11517_));
 sky130_fd_sc_hd__nor2_1 _19099_ (.A(_11516_),
    .B(_11517_),
    .Y(_11518_));
 sky130_fd_sc_hd__xnor2_1 _19100_ (.A(_11512_),
    .B(_11518_),
    .Y(_11519_));
 sky130_fd_sc_hd__nand2_1 _19101_ (.A(_11147_),
    .B(_11161_),
    .Y(_11520_));
 sky130_fd_sc_hd__nor2_1 _19102_ (.A(_11351_),
    .B(_11143_),
    .Y(_11521_));
 sky130_fd_sc_hd__and3_1 _19103_ (.A(_11164_),
    .B(_11145_),
    .C(_11521_),
    .X(_11522_));
 sky130_fd_sc_hd__a21oi_1 _19104_ (.A1(_11164_),
    .A2(_11145_),
    .B1(_11521_),
    .Y(_11523_));
 sky130_fd_sc_hd__nor3_1 _19105_ (.A(_11520_),
    .B(_11522_),
    .C(_11523_),
    .Y(_11524_));
 sky130_fd_sc_hd__o21a_1 _19106_ (.A1(_11522_),
    .A2(_11523_),
    .B1(_11520_),
    .X(_11525_));
 sky130_fd_sc_hd__nor2_1 _19107_ (.A(_11524_),
    .B(_11525_),
    .Y(_11526_));
 sky130_fd_sc_hd__nor2_1 _19108_ (.A(_11480_),
    .B(_11482_),
    .Y(_11527_));
 sky130_fd_sc_hd__xnor2_1 _19109_ (.A(_11526_),
    .B(_11527_),
    .Y(_11528_));
 sky130_fd_sc_hd__nand2_1 _19110_ (.A(_11479_),
    .B(_11528_),
    .Y(_11529_));
 sky130_fd_sc_hd__or2_1 _19111_ (.A(_11479_),
    .B(_11528_),
    .X(_11530_));
 sky130_fd_sc_hd__nand2_1 _19112_ (.A(_11529_),
    .B(_11530_),
    .Y(_11531_));
 sky130_fd_sc_hd__or3_1 _19113_ (.A(_11482_),
    .B(_11484_),
    .C(_11486_),
    .X(_11532_));
 sky130_fd_sc_hd__a21bo_1 _19114_ (.A1(_11479_),
    .A2(_11487_),
    .B1_N(_11532_),
    .X(_11533_));
 sky130_fd_sc_hd__xor2_1 _19115_ (.A(_11531_),
    .B(_11533_),
    .X(_11534_));
 sky130_fd_sc_hd__xor2_1 _19116_ (.A(_11519_),
    .B(_11534_),
    .X(_11535_));
 sky130_fd_sc_hd__or2b_1 _19117_ (.A(_11511_),
    .B_N(_11535_),
    .X(_11536_));
 sky130_fd_sc_hd__or2b_1 _19118_ (.A(_11535_),
    .B_N(_11511_),
    .X(_11537_));
 sky130_fd_sc_hd__nand2_1 _19119_ (.A(_11536_),
    .B(_11537_),
    .Y(_11538_));
 sky130_fd_sc_hd__xnor2_1 _19120_ (.A(_11509_),
    .B(_11538_),
    .Y(_11539_));
 sky130_fd_sc_hd__a21oi_1 _19121_ (.A1(_11506_),
    .A2(_11507_),
    .B1(_11539_),
    .Y(_11540_));
 sky130_fd_sc_hd__and3_1 _19122_ (.A(_11506_),
    .B(_11507_),
    .C(_11539_),
    .X(_11541_));
 sky130_fd_sc_hd__nor2_1 _19123_ (.A(_11540_),
    .B(_11541_),
    .Y(_11542_));
 sky130_fd_sc_hd__xnor2_1 _19124_ (.A(_11498_),
    .B(_11542_),
    .Y(_11543_));
 sky130_fd_sc_hd__nand2_1 _19125_ (.A(_11505_),
    .B(_11543_),
    .Y(_11544_));
 sky130_fd_sc_hd__or2_1 _19126_ (.A(_11505_),
    .B(_11543_),
    .X(_11545_));
 sky130_fd_sc_hd__and2_1 _19127_ (.A(_11544_),
    .B(_11545_),
    .X(_11546_));
 sky130_fd_sc_hd__or2_1 _19128_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[12] ),
    .B(_10639_),
    .X(_11547_));
 sky130_fd_sc_hd__o211a_1 _19129_ (.A1(_11177_),
    .A2(_11546_),
    .B1(_11547_),
    .C1(_11160_),
    .X(_00703_));
 sky130_fd_sc_hd__or3_1 _19130_ (.A(_11498_),
    .B(_11540_),
    .C(_11541_),
    .X(_11548_));
 sky130_fd_sc_hd__a21o_1 _19131_ (.A1(_11506_),
    .A2(_11507_),
    .B1(_11539_),
    .X(_11549_));
 sky130_fd_sc_hd__a21o_1 _19132_ (.A1(_11512_),
    .A2(_11518_),
    .B1(_11516_),
    .X(_11550_));
 sky130_fd_sc_hd__a21o_1 _19133_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[12] ),
    .A2(_11469_),
    .B1(_11387_),
    .X(_11551_));
 sky130_fd_sc_hd__xnor2_1 _19134_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[13] ),
    .B(_11469_),
    .Y(_11552_));
 sky130_fd_sc_hd__nor2_1 _19135_ (.A(_11514_),
    .B(_11552_),
    .Y(_11553_));
 sky130_fd_sc_hd__and2_1 _19136_ (.A(_11514_),
    .B(_11552_),
    .X(_11554_));
 sky130_fd_sc_hd__nor2_1 _19137_ (.A(_11553_),
    .B(_11554_),
    .Y(_11555_));
 sky130_fd_sc_hd__xnor2_2 _19138_ (.A(_11551_),
    .B(_11555_),
    .Y(_11556_));
 sky130_fd_sc_hd__or3_1 _19139_ (.A(_11524_),
    .B(_11525_),
    .C(_11527_),
    .X(_11557_));
 sky130_fd_sc_hd__nand2_1 _19140_ (.A(\top_inst.grid_inst.data_path_wires[13][7] ),
    .B(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[6] ),
    .Y(_11558_));
 sky130_fd_sc_hd__or3_1 _19141_ (.A(_11351_),
    .B(\top_inst.grid_inst.data_path_wires[13][6] ),
    .C(_11558_),
    .X(_11559_));
 sky130_fd_sc_hd__o21ai_1 _19142_ (.A1(_11351_),
    .A2(\top_inst.grid_inst.data_path_wires[13][6] ),
    .B1(_11558_),
    .Y(_11560_));
 sky130_fd_sc_hd__and2_1 _19143_ (.A(_11559_),
    .B(_11560_),
    .X(_11561_));
 sky130_fd_sc_hd__xnor2_1 _19144_ (.A(_11520_),
    .B(_11561_),
    .Y(_11562_));
 sky130_fd_sc_hd__o21ai_1 _19145_ (.A1(_11522_),
    .A2(_11524_),
    .B1(_11562_),
    .Y(_11563_));
 sky130_fd_sc_hd__or3_1 _19146_ (.A(_11522_),
    .B(_11524_),
    .C(_11562_),
    .X(_11564_));
 sky130_fd_sc_hd__and2_1 _19147_ (.A(_11563_),
    .B(_11564_),
    .X(_11565_));
 sky130_fd_sc_hd__nand2_1 _19148_ (.A(_11479_),
    .B(_11565_),
    .Y(_11566_));
 sky130_fd_sc_hd__or2_1 _19149_ (.A(_11479_),
    .B(_11565_),
    .X(_11567_));
 sky130_fd_sc_hd__nand2_1 _19150_ (.A(_11566_),
    .B(_11567_),
    .Y(_11568_));
 sky130_fd_sc_hd__a21o_1 _19151_ (.A1(_11557_),
    .A2(_11529_),
    .B1(_11568_),
    .X(_11569_));
 sky130_fd_sc_hd__nand3_1 _19152_ (.A(_11557_),
    .B(_11529_),
    .C(_11568_),
    .Y(_11570_));
 sky130_fd_sc_hd__nand2_1 _19153_ (.A(_11569_),
    .B(_11570_),
    .Y(_11571_));
 sky130_fd_sc_hd__xor2_2 _19154_ (.A(_11556_),
    .B(_11571_),
    .X(_11572_));
 sky130_fd_sc_hd__or2b_1 _19155_ (.A(_11531_),
    .B_N(_11533_),
    .X(_11573_));
 sky130_fd_sc_hd__o21a_1 _19156_ (.A1(_11519_),
    .A2(_11534_),
    .B1(_11573_),
    .X(_11574_));
 sky130_fd_sc_hd__xor2_1 _19157_ (.A(_11572_),
    .B(_11574_),
    .X(_11575_));
 sky130_fd_sc_hd__xor2_1 _19158_ (.A(_11550_),
    .B(_11575_),
    .X(_11576_));
 sky130_fd_sc_hd__o21a_1 _19159_ (.A1(_11509_),
    .A2(_11538_),
    .B1(_11536_),
    .X(_11577_));
 sky130_fd_sc_hd__or2_1 _19160_ (.A(_11576_),
    .B(_11577_),
    .X(_11578_));
 sky130_fd_sc_hd__nand2_1 _19161_ (.A(_11576_),
    .B(_11577_),
    .Y(_11579_));
 sky130_fd_sc_hd__and2_1 _19162_ (.A(_11578_),
    .B(_11579_),
    .X(_11580_));
 sky130_fd_sc_hd__xnor2_1 _19163_ (.A(_11549_),
    .B(_11580_),
    .Y(_11581_));
 sky130_fd_sc_hd__a21oi_1 _19164_ (.A1(_11548_),
    .A2(_11544_),
    .B1(_11581_),
    .Y(_11582_));
 sky130_fd_sc_hd__a31o_1 _19165_ (.A1(_11548_),
    .A2(_11544_),
    .A3(_11581_),
    .B1(_10957_),
    .X(_11583_));
 sky130_fd_sc_hd__o221a_1 _19166_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[13] ),
    .A2(_10364_),
    .B1(_11582_),
    .B2(_11583_),
    .C1(_11228_),
    .X(_00704_));
 sky130_fd_sc_hd__nand2_1 _19167_ (.A(_11549_),
    .B(_11548_),
    .Y(_11584_));
 sky130_fd_sc_hd__a32o_1 _19168_ (.A1(_11505_),
    .A2(_11543_),
    .A3(_11581_),
    .B1(_11584_),
    .B2(_11580_),
    .X(_11585_));
 sky130_fd_sc_hd__a21o_1 _19169_ (.A1(_11551_),
    .A2(_11555_),
    .B1(_11553_),
    .X(_11586_));
 sky130_fd_sc_hd__inv_2 _19170_ (.A(_11586_),
    .Y(_11587_));
 sky130_fd_sc_hd__o21a_1 _19171_ (.A1(_11556_),
    .A2(_11571_),
    .B1(_11569_),
    .X(_11588_));
 sky130_fd_sc_hd__a21o_1 _19172_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[13] ),
    .A2(_11469_),
    .B1(_11387_),
    .X(_11589_));
 sky130_fd_sc_hd__and2_1 _19173_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[14] ),
    .B(_11469_),
    .X(_11590_));
 sky130_fd_sc_hd__nor2_1 _19174_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[14] ),
    .B(_11469_),
    .Y(_11591_));
 sky130_fd_sc_hd__or2_1 _19175_ (.A(_11590_),
    .B(_11591_),
    .X(_11592_));
 sky130_fd_sc_hd__xor2_1 _19176_ (.A(_11514_),
    .B(_11592_),
    .X(_11593_));
 sky130_fd_sc_hd__nand2_1 _19177_ (.A(_11589_),
    .B(_11593_),
    .Y(_11594_));
 sky130_fd_sc_hd__or2_1 _19178_ (.A(_11589_),
    .B(_11593_),
    .X(_11595_));
 sky130_fd_sc_hd__nand2_1 _19179_ (.A(_11594_),
    .B(_11595_),
    .Y(_11596_));
 sky130_fd_sc_hd__o211a_1 _19180_ (.A1(_11351_),
    .A2(_11147_),
    .B1(_11520_),
    .C1(_11558_),
    .X(_11597_));
 sky130_fd_sc_hd__and2_1 _19181_ (.A(_11147_),
    .B(_11161_),
    .X(_11598_));
 sky130_fd_sc_hd__nand2_1 _19182_ (.A(_11598_),
    .B(_11561_),
    .Y(_11599_));
 sky130_fd_sc_hd__a22oi_2 _19183_ (.A1(_11164_),
    .A2(_11598_),
    .B1(_11559_),
    .B2(_11599_),
    .Y(_11600_));
 sky130_fd_sc_hd__nor2_1 _19184_ (.A(_11597_),
    .B(_11600_),
    .Y(_11601_));
 sky130_fd_sc_hd__xnor2_1 _19185_ (.A(_11479_),
    .B(_11601_),
    .Y(_11602_));
 sky130_fd_sc_hd__a21oi_1 _19186_ (.A1(_11563_),
    .A2(_11566_),
    .B1(_11602_),
    .Y(_11603_));
 sky130_fd_sc_hd__and3_1 _19187_ (.A(_11563_),
    .B(_11566_),
    .C(_11602_),
    .X(_11604_));
 sky130_fd_sc_hd__nor2_1 _19188_ (.A(_11603_),
    .B(_11604_),
    .Y(_11605_));
 sky130_fd_sc_hd__xnor2_1 _19189_ (.A(_11596_),
    .B(_11605_),
    .Y(_11606_));
 sky130_fd_sc_hd__or2b_1 _19190_ (.A(_11588_),
    .B_N(_11606_),
    .X(_11607_));
 sky130_fd_sc_hd__or2b_1 _19191_ (.A(_11606_),
    .B_N(_11588_),
    .X(_11608_));
 sky130_fd_sc_hd__nand2_1 _19192_ (.A(_11607_),
    .B(_11608_),
    .Y(_11609_));
 sky130_fd_sc_hd__xnor2_2 _19193_ (.A(_11587_),
    .B(_11609_),
    .Y(_11610_));
 sky130_fd_sc_hd__inv_2 _19194_ (.A(_11574_),
    .Y(_11611_));
 sky130_fd_sc_hd__and2b_1 _19195_ (.A_N(_11575_),
    .B(_11550_),
    .X(_11612_));
 sky130_fd_sc_hd__a21oi_2 _19196_ (.A1(_11572_),
    .A2(_11611_),
    .B1(_11612_),
    .Y(_11613_));
 sky130_fd_sc_hd__xor2_2 _19197_ (.A(_11610_),
    .B(_11613_),
    .X(_11614_));
 sky130_fd_sc_hd__xnor2_2 _19198_ (.A(_11578_),
    .B(_11614_),
    .Y(_11615_));
 sky130_fd_sc_hd__xor2_1 _19199_ (.A(_11585_),
    .B(_11615_),
    .X(_11616_));
 sky130_fd_sc_hd__or2_1 _19200_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[14] ),
    .B(_10639_),
    .X(_11617_));
 sky130_fd_sc_hd__o211a_1 _19201_ (.A1(_11177_),
    .A2(_11616_),
    .B1(_11617_),
    .C1(_11160_),
    .X(_00705_));
 sky130_fd_sc_hd__or2b_1 _19202_ (.A(_11578_),
    .B_N(_11614_),
    .X(_11618_));
 sky130_fd_sc_hd__a21boi_1 _19203_ (.A1(_11585_),
    .A2(_11615_),
    .B1_N(_11618_),
    .Y(_11619_));
 sky130_fd_sc_hd__or2_1 _19204_ (.A(_11610_),
    .B(_11613_),
    .X(_11620_));
 sky130_fd_sc_hd__o21ai_1 _19205_ (.A1(_11514_),
    .A2(_11592_),
    .B1(_11594_),
    .Y(_11621_));
 sky130_fd_sc_hd__nor2_1 _19206_ (.A(_11479_),
    .B(_11601_),
    .Y(_11622_));
 sky130_fd_sc_hd__xnor2_1 _19207_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[15] ),
    .B(_11469_),
    .Y(_11623_));
 sky130_fd_sc_hd__nor2_1 _19208_ (.A(_11514_),
    .B(_11623_),
    .Y(_11624_));
 sky130_fd_sc_hd__and2_1 _19209_ (.A(_11514_),
    .B(_11623_),
    .X(_11625_));
 sky130_fd_sc_hd__nor2_1 _19210_ (.A(_11624_),
    .B(_11625_),
    .Y(_11626_));
 sky130_fd_sc_hd__o21a_1 _19211_ (.A1(_11387_),
    .A2(_11590_),
    .B1(_11626_),
    .X(_11627_));
 sky130_fd_sc_hd__nor3_1 _19212_ (.A(_11387_),
    .B(_11590_),
    .C(_11626_),
    .Y(_11628_));
 sky130_fd_sc_hd__or2_1 _19213_ (.A(_11627_),
    .B(_11628_),
    .X(_11629_));
 sky130_fd_sc_hd__xor2_2 _19214_ (.A(_11622_),
    .B(_11629_),
    .X(_11630_));
 sky130_fd_sc_hd__a31o_1 _19215_ (.A1(_11594_),
    .A2(_11595_),
    .A3(_11605_),
    .B1(_11603_),
    .X(_11631_));
 sky130_fd_sc_hd__xnor2_1 _19216_ (.A(_11630_),
    .B(_11631_),
    .Y(_11632_));
 sky130_fd_sc_hd__xor2_1 _19217_ (.A(_11621_),
    .B(_11632_),
    .X(_11633_));
 sky130_fd_sc_hd__o21a_1 _19218_ (.A1(_11587_),
    .A2(_11609_),
    .B1(_11607_),
    .X(_11634_));
 sky130_fd_sc_hd__or2_1 _19219_ (.A(_11633_),
    .B(_11634_),
    .X(_11635_));
 sky130_fd_sc_hd__nand2_1 _19220_ (.A(_11633_),
    .B(_11634_),
    .Y(_11636_));
 sky130_fd_sc_hd__and2_1 _19221_ (.A(_11635_),
    .B(_11636_),
    .X(_11637_));
 sky130_fd_sc_hd__xnor2_1 _19222_ (.A(_11620_),
    .B(_11637_),
    .Y(_11638_));
 sky130_fd_sc_hd__nor2_1 _19223_ (.A(_11619_),
    .B(_11638_),
    .Y(_11639_));
 sky130_fd_sc_hd__a2111o_1 _19224_ (.A1(_11619_),
    .A2(_11638_),
    .B1(_11639_),
    .C1(_05309_),
    .D1(_04861_),
    .X(_11640_));
 sky130_fd_sc_hd__buf_4 _19225_ (.A(_10447_),
    .X(_11641_));
 sky130_fd_sc_hd__o211a_1 _19226_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[15] ),
    .A2(_10616_),
    .B1(_11640_),
    .C1(_11641_),
    .X(_00706_));
 sky130_fd_sc_hd__nand2_1 _19227_ (.A(_11620_),
    .B(_11618_),
    .Y(_11642_));
 sky130_fd_sc_hd__a32o_1 _19228_ (.A1(_11585_),
    .A2(_11615_),
    .A3(_11638_),
    .B1(_11642_),
    .B2(_11637_),
    .X(_11643_));
 sky130_fd_sc_hd__inv_2 _19229_ (.A(_11479_),
    .Y(_11644_));
 sky130_fd_sc_hd__o2bb2a_1 _19230_ (.A1_N(_11644_),
    .A2_N(_11600_),
    .B1(_11622_),
    .B2(_11629_),
    .X(_11645_));
 sky130_fd_sc_hd__nand2_1 _19231_ (.A(_11644_),
    .B(_11597_),
    .Y(_11646_));
 sky130_fd_sc_hd__a21o_1 _19232_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[15] ),
    .A2(_11469_),
    .B1(_11387_),
    .X(_11647_));
 sky130_fd_sc_hd__xnor2_2 _19233_ (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[16] ),
    .B(_11469_),
    .Y(_11648_));
 sky130_fd_sc_hd__xor2_1 _19234_ (.A(_11514_),
    .B(_11648_),
    .X(_11649_));
 sky130_fd_sc_hd__xnor2_1 _19235_ (.A(_11647_),
    .B(_11649_),
    .Y(_11650_));
 sky130_fd_sc_hd__xor2_1 _19236_ (.A(_11646_),
    .B(_11650_),
    .X(_11651_));
 sky130_fd_sc_hd__xor2_1 _19237_ (.A(_11645_),
    .B(_11651_),
    .X(_11652_));
 sky130_fd_sc_hd__o21ai_1 _19238_ (.A1(_11624_),
    .A2(_11627_),
    .B1(_11652_),
    .Y(_11653_));
 sky130_fd_sc_hd__or3_1 _19239_ (.A(_11624_),
    .B(_11627_),
    .C(_11652_),
    .X(_11654_));
 sky130_fd_sc_hd__nand2_1 _19240_ (.A(_11653_),
    .B(_11654_),
    .Y(_11655_));
 sky130_fd_sc_hd__and2b_1 _19241_ (.A_N(_11632_),
    .B(_11621_),
    .X(_11656_));
 sky130_fd_sc_hd__a21oi_1 _19242_ (.A1(_11630_),
    .A2(_11631_),
    .B1(_11656_),
    .Y(_11657_));
 sky130_fd_sc_hd__xor2_1 _19243_ (.A(_11655_),
    .B(_11657_),
    .X(_11658_));
 sky130_fd_sc_hd__xnor2_1 _19244_ (.A(_11635_),
    .B(_11658_),
    .Y(_11659_));
 sky130_fd_sc_hd__xor2_1 _19245_ (.A(_11643_),
    .B(_11659_),
    .X(_11660_));
 sky130_fd_sc_hd__or2_1 _19246_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[16] ),
    .B(_10639_),
    .X(_11661_));
 sky130_fd_sc_hd__o211a_1 _19247_ (.A1(_11177_),
    .A2(_11660_),
    .B1(_11661_),
    .C1(_11641_),
    .X(_00707_));
 sky130_fd_sc_hd__clkbuf_4 _19248_ (.A(_05313_),
    .X(_11662_));
 sky130_fd_sc_hd__nor2_1 _19249_ (.A(_11655_),
    .B(_11657_),
    .Y(_11663_));
 sky130_fd_sc_hd__o21a_1 _19250_ (.A1(_11645_),
    .A2(_11651_),
    .B1(_11653_),
    .X(_11664_));
 sky130_fd_sc_hd__a21o_1 _19251_ (.A1(_11514_),
    .A2(_11648_),
    .B1(_11647_),
    .X(_11665_));
 sky130_fd_sc_hd__o21a_1 _19252_ (.A1(_11514_),
    .A2(_11648_),
    .B1(_11665_),
    .X(_11666_));
 sky130_fd_sc_hd__nand2_1 _19253_ (.A(_11646_),
    .B(_11650_),
    .Y(_11667_));
 sky130_fd_sc_hd__o21ba_1 _19254_ (.A1(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[16] ),
    .A2(_11387_),
    .B1_N(_11338_),
    .X(_11668_));
 sky130_fd_sc_hd__xnor2_1 _19255_ (.A(_11667_),
    .B(_11668_),
    .Y(_11669_));
 sky130_fd_sc_hd__xnor2_1 _19256_ (.A(_11666_),
    .B(_11669_),
    .Y(_11670_));
 sky130_fd_sc_hd__xnor2_1 _19257_ (.A(_11664_),
    .B(_11670_),
    .Y(_11671_));
 sky130_fd_sc_hd__xnor2_1 _19258_ (.A(_11663_),
    .B(_11671_),
    .Y(_11672_));
 sky130_fd_sc_hd__and2b_1 _19259_ (.A_N(_11635_),
    .B(_11658_),
    .X(_11673_));
 sky130_fd_sc_hd__a211o_1 _19260_ (.A1(_11643_),
    .A2(_11659_),
    .B1(_11672_),
    .C1(_11673_),
    .X(_11674_));
 sky130_fd_sc_hd__a21oi_4 _19261_ (.A1(_05787_),
    .A2(_11674_),
    .B1(_04867_),
    .Y(_11675_));
 sky130_fd_sc_hd__o21a_1 _19262_ (.A1(net963),
    .A2(_11662_),
    .B1(_11675_),
    .X(_00708_));
 sky130_fd_sc_hd__o21a_1 _19263_ (.A1(net957),
    .A2(_11662_),
    .B1(_11675_),
    .X(_00709_));
 sky130_fd_sc_hd__o21a_1 _19264_ (.A1(net959),
    .A2(_11662_),
    .B1(_11675_),
    .X(_00710_));
 sky130_fd_sc_hd__o21a_1 _19265_ (.A1(net960),
    .A2(_11662_),
    .B1(_11675_),
    .X(_00711_));
 sky130_fd_sc_hd__o21a_1 _19266_ (.A1(net1018),
    .A2(_11662_),
    .B1(_11675_),
    .X(_00712_));
 sky130_fd_sc_hd__o21a_1 _19267_ (.A1(net962),
    .A2(_11662_),
    .B1(_11675_),
    .X(_00713_));
 sky130_fd_sc_hd__o21a_1 _19268_ (.A1(net985),
    .A2(_11662_),
    .B1(_11675_),
    .X(_00714_));
 sky130_fd_sc_hd__o21a_1 _19269_ (.A1(net1057),
    .A2(_11662_),
    .B1(_11675_),
    .X(_00715_));
 sky130_fd_sc_hd__o21a_1 _19270_ (.A1(net1032),
    .A2(_11662_),
    .B1(_11675_),
    .X(_00716_));
 sky130_fd_sc_hd__o21a_1 _19271_ (.A1(net748),
    .A2(_11662_),
    .B1(_11675_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_2 _19272_ (.A0(\top_inst.skew_buff_inst.row[3].output_reg[0] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[24] ),
    .S(net205),
    .X(_11676_));
 sky130_fd_sc_hd__buf_2 _19273_ (.A(net245),
    .X(_11677_));
 sky130_fd_sc_hd__buf_2 _19274_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[0] ),
    .X(_11678_));
 sky130_fd_sc_hd__clkbuf_4 _19275_ (.A(_11678_),
    .X(_11679_));
 sky130_fd_sc_hd__or2_1 _19276_ (.A(_11679_),
    .B(_11150_),
    .X(_11680_));
 sky130_fd_sc_hd__o211a_1 _19277_ (.A1(_09185_),
    .A2(_11677_),
    .B1(_11680_),
    .C1(_11641_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_4 _19278_ (.A0(\top_inst.skew_buff_inst.row[3].output_reg[1] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[25] ),
    .S(net188),
    .X(_11681_));
 sky130_fd_sc_hd__buf_2 _19279_ (.A(net190),
    .X(_11682_));
 sky130_fd_sc_hd__clkbuf_4 _19280_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[1] ),
    .X(_11683_));
 sky130_fd_sc_hd__clkbuf_4 _19281_ (.A(_11683_),
    .X(_11684_));
 sky130_fd_sc_hd__or2_1 _19282_ (.A(_11684_),
    .B(_11150_),
    .X(_11685_));
 sky130_fd_sc_hd__o211a_1 _19283_ (.A1(_09185_),
    .A2(_11682_),
    .B1(_11685_),
    .C1(_11641_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_4 _19284_ (.A0(\top_inst.skew_buff_inst.row[3].output_reg[2] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[26] ),
    .S(net188),
    .X(_11686_));
 sky130_fd_sc_hd__buf_6 _19285_ (.A(net247),
    .X(_11687_));
 sky130_fd_sc_hd__clkbuf_4 _19286_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[2] ),
    .X(_11688_));
 sky130_fd_sc_hd__clkbuf_4 _19287_ (.A(_05772_),
    .X(_11689_));
 sky130_fd_sc_hd__or2_1 _19288_ (.A(_11688_),
    .B(_11689_),
    .X(_11690_));
 sky130_fd_sc_hd__o211a_1 _19289_ (.A1(_09185_),
    .A2(_11687_),
    .B1(_11690_),
    .C1(_11641_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_4 _19290_ (.A0(\top_inst.skew_buff_inst.row[3].output_reg[3] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[27] ),
    .S(net184),
    .X(_11691_));
 sky130_fd_sc_hd__buf_4 _19291_ (.A(net240),
    .X(_11692_));
 sky130_fd_sc_hd__clkbuf_4 _19292_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[3] ),
    .X(_11693_));
 sky130_fd_sc_hd__or2_1 _19293_ (.A(_11693_),
    .B(_11689_),
    .X(_11694_));
 sky130_fd_sc_hd__o211a_1 _19294_ (.A1(_09185_),
    .A2(_11692_),
    .B1(_11694_),
    .C1(_11641_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_4 _19295_ (.A0(\top_inst.skew_buff_inst.row[3].output_reg[4] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[28] ),
    .S(net34),
    .X(_11695_));
 sky130_fd_sc_hd__clkbuf_4 _19296_ (.A(_11695_),
    .X(_11696_));
 sky130_fd_sc_hd__clkbuf_4 _19297_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[4] ),
    .X(_11697_));
 sky130_fd_sc_hd__or2_1 _19298_ (.A(_11697_),
    .B(_11689_),
    .X(_11698_));
 sky130_fd_sc_hd__o211a_1 _19299_ (.A1(_05755_),
    .A2(_11696_),
    .B1(_11698_),
    .C1(_11641_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_4 _19300_ (.A0(\top_inst.skew_buff_inst.row[3].output_reg[5] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[29] ),
    .S(net188),
    .X(_11699_));
 sky130_fd_sc_hd__clkbuf_4 _19301_ (.A(net193),
    .X(_11700_));
 sky130_fd_sc_hd__buf_2 _19302_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[5] ),
    .X(_11701_));
 sky130_fd_sc_hd__or2_1 _19303_ (.A(_11701_),
    .B(_11689_),
    .X(_11702_));
 sky130_fd_sc_hd__o211a_1 _19304_ (.A1(_05755_),
    .A2(_11700_),
    .B1(_11702_),
    .C1(_11641_),
    .X(_00723_));
 sky130_fd_sc_hd__buf_2 _19305_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[6] ),
    .X(_11703_));
 sky130_fd_sc_hd__mux2_4 _19306_ (.A0(\top_inst.skew_buff_inst.row[3].output_reg[6] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[30] ),
    .S(net188),
    .X(_11704_));
 sky130_fd_sc_hd__buf_2 _19307_ (.A(_11704_),
    .X(_11705_));
 sky130_fd_sc_hd__or2_1 _19308_ (.A(_05269_),
    .B(_11705_),
    .X(_11706_));
 sky130_fd_sc_hd__o211a_1 _19309_ (.A1(_11703_),
    .A2(_05276_),
    .B1(_11706_),
    .C1(_11641_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_2 _19310_ (.A0(\top_inst.skew_buff_inst.row[3].output_reg[7] ),
    .A1(\top_inst.axis_in_inst.inbuf_bus[31] ),
    .S(net34),
    .X(_11707_));
 sky130_fd_sc_hd__clkbuf_4 _19311_ (.A(_11707_),
    .X(_11708_));
 sky130_fd_sc_hd__clkbuf_4 _19312_ (.A(_11708_),
    .X(_11709_));
 sky130_fd_sc_hd__or2_1 _19313_ (.A(_05269_),
    .B(_11709_),
    .X(_11710_));
 sky130_fd_sc_hd__o211a_1 _19314_ (.A1(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[7] ),
    .A2(_05276_),
    .B1(_11710_),
    .C1(_11641_),
    .X(_00725_));
 sky130_fd_sc_hd__a21oi_1 _19315_ (.A1(_11679_),
    .A2(_11677_),
    .B1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[0] ),
    .Y(_11711_));
 sky130_fd_sc_hd__and3_1 _19316_ (.A(_11679_),
    .B(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[0] ),
    .C(_11677_),
    .X(_11712_));
 sky130_fd_sc_hd__o21ai_2 _19317_ (.A1(_11711_),
    .A2(_11712_),
    .B1(_08181_),
    .Y(_11713_));
 sky130_fd_sc_hd__buf_2 _19318_ (.A(_10447_),
    .X(_11714_));
 sky130_fd_sc_hd__o211a_1 _19319_ (.A1(net917),
    .A2(_10616_),
    .B1(_11713_),
    .C1(_11714_),
    .X(_00726_));
 sky130_fd_sc_hd__a22o_1 _19320_ (.A1(_11684_),
    .A2(_11677_),
    .B1(_11682_),
    .B2(_11679_),
    .X(_11715_));
 sky130_fd_sc_hd__nand4_1 _19321_ (.A(_11684_),
    .B(_11679_),
    .C(_11677_),
    .D(_11682_),
    .Y(_11716_));
 sky130_fd_sc_hd__and3_1 _19322_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[1] ),
    .B(_11715_),
    .C(_11716_),
    .X(_11717_));
 sky130_fd_sc_hd__a21oi_1 _19323_ (.A1(_11715_),
    .A2(_11716_),
    .B1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[1] ),
    .Y(_11718_));
 sky130_fd_sc_hd__o21ba_1 _19324_ (.A1(_11717_),
    .A2(_11718_),
    .B1_N(_11712_),
    .X(_11719_));
 sky130_fd_sc_hd__nor3b_1 _19325_ (.A(_11717_),
    .B(_11718_),
    .C_N(_11712_),
    .Y(_11720_));
 sky130_fd_sc_hd__o21ai_2 _19326_ (.A1(_11719_),
    .A2(_11720_),
    .B1(_08181_),
    .Y(_11721_));
 sky130_fd_sc_hd__o211a_1 _19327_ (.A1(net932),
    .A2(_10616_),
    .B1(_11721_),
    .C1(_11714_),
    .X(_00727_));
 sky130_fd_sc_hd__clkbuf_4 _19328_ (.A(_04873_),
    .X(_11722_));
 sky130_fd_sc_hd__buf_6 _19329_ (.A(_05326_),
    .X(_11723_));
 sky130_fd_sc_hd__nand2_1 _19330_ (.A(_11688_),
    .B(_11677_),
    .Y(_11724_));
 sky130_fd_sc_hd__a22o_1 _19331_ (.A1(_11684_),
    .A2(_11682_),
    .B1(_11687_),
    .B2(_11679_),
    .X(_11725_));
 sky130_fd_sc_hd__nand4_2 _19332_ (.A(_11684_),
    .B(_11679_),
    .C(_11682_),
    .D(_11687_),
    .Y(_11726_));
 sky130_fd_sc_hd__nand3_1 _19333_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[2] ),
    .B(_11725_),
    .C(_11726_),
    .Y(_11727_));
 sky130_fd_sc_hd__a21o_1 _19334_ (.A1(_11725_),
    .A2(_11726_),
    .B1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[2] ),
    .X(_11728_));
 sky130_fd_sc_hd__nand2_1 _19335_ (.A(_11727_),
    .B(_11728_),
    .Y(_11729_));
 sky130_fd_sc_hd__a21boi_1 _19336_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[1] ),
    .A2(_11715_),
    .B1_N(_11716_),
    .Y(_11730_));
 sky130_fd_sc_hd__xnor2_1 _19337_ (.A(_11729_),
    .B(_11730_),
    .Y(_11731_));
 sky130_fd_sc_hd__xor2_1 _19338_ (.A(_11724_),
    .B(_11731_),
    .X(_11732_));
 sky130_fd_sc_hd__nand2_1 _19339_ (.A(net172),
    .B(_11732_),
    .Y(_01178_));
 sky130_fd_sc_hd__o21a_1 _19340_ (.A1(net172),
    .A2(_11732_),
    .B1(_10831_),
    .X(_01179_));
 sky130_fd_sc_hd__a22o_1 _19341_ (.A1(\top_inst.deskew_buff_inst.col_input[2] ),
    .A2(_11723_),
    .B1(_01178_),
    .B2(_01179_),
    .X(_01180_));
 sky130_fd_sc_hd__and2_1 _19342_ (.A(_11722_),
    .B(_01180_),
    .X(_01181_));
 sky130_fd_sc_hd__clkbuf_1 _19343_ (.A(_01181_),
    .X(_00728_));
 sky130_fd_sc_hd__or2_1 _19344_ (.A(_11729_),
    .B(_11730_),
    .X(_01182_));
 sky130_fd_sc_hd__or2_1 _19345_ (.A(_11724_),
    .B(_11731_),
    .X(_01183_));
 sky130_fd_sc_hd__a22o_1 _19346_ (.A1(_11693_),
    .A2(_11677_),
    .B1(_11682_),
    .B2(_11688_),
    .X(_01184_));
 sky130_fd_sc_hd__nand4_1 _19347_ (.A(_11693_),
    .B(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[2] ),
    .C(net243),
    .D(_11682_),
    .Y(_01185_));
 sky130_fd_sc_hd__and2_1 _19348_ (.A(_01184_),
    .B(_01185_),
    .X(_01186_));
 sky130_fd_sc_hd__a22o_1 _19349_ (.A1(_11683_),
    .A2(_11687_),
    .B1(_11692_),
    .B2(_11678_),
    .X(_01187_));
 sky130_fd_sc_hd__nand4_1 _19350_ (.A(_11684_),
    .B(_11679_),
    .C(_11687_),
    .D(_11692_),
    .Y(_01188_));
 sky130_fd_sc_hd__and3_1 _19351_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[3] ),
    .B(_01187_),
    .C(_01188_),
    .X(_01189_));
 sky130_fd_sc_hd__a21oi_1 _19352_ (.A1(_01187_),
    .A2(_01188_),
    .B1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[3] ),
    .Y(_01190_));
 sky130_fd_sc_hd__a211oi_1 _19353_ (.A1(_11726_),
    .A2(_11727_),
    .B1(_01189_),
    .C1(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__o211ai_1 _19354_ (.A1(_01189_),
    .A2(_01190_),
    .B1(_11726_),
    .C1(_11727_),
    .Y(_01192_));
 sky130_fd_sc_hd__or2b_1 _19355_ (.A(_01191_),
    .B_N(_01192_),
    .X(_01193_));
 sky130_fd_sc_hd__xor2_1 _19356_ (.A(_01186_),
    .B(_01193_),
    .X(_01194_));
 sky130_fd_sc_hd__a21oi_2 _19357_ (.A1(_01182_),
    .A2(_01183_),
    .B1(_01194_),
    .Y(_01195_));
 sky130_fd_sc_hd__and3_1 _19358_ (.A(_01182_),
    .B(_01183_),
    .C(_01194_),
    .X(_01196_));
 sky130_fd_sc_hd__or3_1 _19359_ (.A(_01178_),
    .B(_01195_),
    .C(_01196_),
    .X(_01197_));
 sky130_fd_sc_hd__o21ai_1 _19360_ (.A1(_01195_),
    .A2(_01196_),
    .B1(_01178_),
    .Y(_01198_));
 sky130_fd_sc_hd__and2_1 _19361_ (.A(\top_inst.deskew_buff_inst.col_input[3] ),
    .B(_05730_),
    .X(_01199_));
 sky130_fd_sc_hd__a31o_1 _19362_ (.A1(_05887_),
    .A2(_01197_),
    .A3(_01198_),
    .B1(_01199_),
    .X(_01200_));
 sky130_fd_sc_hd__and2_1 _19363_ (.A(_11722_),
    .B(_01200_),
    .X(_01201_));
 sky130_fd_sc_hd__clkbuf_1 _19364_ (.A(_01201_),
    .X(_00729_));
 sky130_fd_sc_hd__buf_4 _19365_ (.A(_06168_),
    .X(_01202_));
 sky130_fd_sc_hd__a22o_1 _19366_ (.A1(_11683_),
    .A2(net233),
    .B1(_11695_),
    .B2(_11678_),
    .X(_01203_));
 sky130_fd_sc_hd__nand4_1 _19367_ (.A(_11683_),
    .B(_11678_),
    .C(net234),
    .D(_11696_),
    .Y(_01204_));
 sky130_fd_sc_hd__and3_1 _19368_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[4] ),
    .B(_01203_),
    .C(_01204_),
    .X(_01205_));
 sky130_fd_sc_hd__a21oi_1 _19369_ (.A1(_01203_),
    .A2(_01204_),
    .B1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[4] ),
    .Y(_01206_));
 sky130_fd_sc_hd__or3_4 _19370_ (.A(_01185_),
    .B(_01205_),
    .C(_01206_),
    .X(_01207_));
 sky130_fd_sc_hd__o21ai_1 _19371_ (.A1(_01205_),
    .A2(_01206_),
    .B1(_01185_),
    .Y(_01208_));
 sky130_fd_sc_hd__a21bo_1 _19372_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[3] ),
    .A2(_01187_),
    .B1_N(_01188_),
    .X(_01209_));
 sky130_fd_sc_hd__nand3_1 _19373_ (.A(_01207_),
    .B(_01208_),
    .C(_01209_),
    .Y(_01210_));
 sky130_fd_sc_hd__a21o_1 _19374_ (.A1(_01207_),
    .A2(_01208_),
    .B1(_01209_),
    .X(_01211_));
 sky130_fd_sc_hd__nand2_1 _19375_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[2] ),
    .B(_11687_),
    .Y(_01212_));
 sky130_fd_sc_hd__nand4_2 _19376_ (.A(_11697_),
    .B(_11693_),
    .C(net243),
    .D(net191),
    .Y(_01213_));
 sky130_fd_sc_hd__a22o_1 _19377_ (.A1(_11697_),
    .A2(net243),
    .B1(net191),
    .B2(_11693_),
    .X(_01214_));
 sky130_fd_sc_hd__nand3b_1 _19378_ (.A_N(_01212_),
    .B(_01213_),
    .C(_01214_),
    .Y(_01215_));
 sky130_fd_sc_hd__a21bo_1 _19379_ (.A1(_01213_),
    .A2(_01214_),
    .B1_N(_01212_),
    .X(_01216_));
 sky130_fd_sc_hd__and2_1 _19380_ (.A(_01215_),
    .B(_01216_),
    .X(_01217_));
 sky130_fd_sc_hd__and3_1 _19381_ (.A(_01210_),
    .B(_01211_),
    .C(_01217_),
    .X(_01218_));
 sky130_fd_sc_hd__a21oi_2 _19382_ (.A1(_01210_),
    .A2(_01211_),
    .B1(_01217_),
    .Y(_01219_));
 sky130_fd_sc_hd__a21o_1 _19383_ (.A1(_01186_),
    .A2(_01192_),
    .B1(_01191_),
    .X(_01220_));
 sky130_fd_sc_hd__or3b_4 _19384_ (.A(_01218_),
    .B(_01219_),
    .C_N(_01220_),
    .X(_01221_));
 sky130_fd_sc_hd__o21bai_2 _19385_ (.A1(_01218_),
    .A2(_01219_),
    .B1_N(_01220_),
    .Y(_01222_));
 sky130_fd_sc_hd__nand2_1 _19386_ (.A(_01221_),
    .B(_01222_),
    .Y(_01223_));
 sky130_fd_sc_hd__or2b_1 _19387_ (.A(_01195_),
    .B_N(_01197_),
    .X(_01224_));
 sky130_fd_sc_hd__nor2_1 _19388_ (.A(_01223_),
    .B(_01224_),
    .Y(_01225_));
 sky130_fd_sc_hd__a21o_1 _19389_ (.A1(_01223_),
    .A2(_01224_),
    .B1(_09292_),
    .X(_01226_));
 sky130_fd_sc_hd__o221a_1 _19390_ (.A1(net355),
    .A2(_01202_),
    .B1(_01225_),
    .B2(_01226_),
    .C1(_11228_),
    .X(_00730_));
 sky130_fd_sc_hd__and2_1 _19391_ (.A(net812),
    .B(_05634_),
    .X(_01227_));
 sky130_fd_sc_hd__nor2_1 _19392_ (.A(_01197_),
    .B(_01223_),
    .Y(_01228_));
 sky130_fd_sc_hd__a21bo_1 _19393_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[4] ),
    .A2(_01203_),
    .B1_N(_01204_),
    .X(_01229_));
 sky130_fd_sc_hd__a22o_1 _19394_ (.A1(_11683_),
    .A2(_11695_),
    .B1(_11700_),
    .B2(_11678_),
    .X(_01230_));
 sky130_fd_sc_hd__nand4_1 _19395_ (.A(_11683_),
    .B(_11678_),
    .C(_11696_),
    .D(_11700_),
    .Y(_01231_));
 sky130_fd_sc_hd__and3_1 _19396_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[5] ),
    .B(_01230_),
    .C(_01231_),
    .X(_01232_));
 sky130_fd_sc_hd__a21oi_1 _19397_ (.A1(_01230_),
    .A2(_01231_),
    .B1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[5] ),
    .Y(_01233_));
 sky130_fd_sc_hd__a211o_1 _19398_ (.A1(_01213_),
    .A2(_01215_),
    .B1(_01232_),
    .C1(_01233_),
    .X(_01234_));
 sky130_fd_sc_hd__o211ai_2 _19399_ (.A1(_01232_),
    .A2(_01233_),
    .B1(_01213_),
    .C1(_01215_),
    .Y(_01235_));
 sky130_fd_sc_hd__nand3_2 _19400_ (.A(_01229_),
    .B(_01234_),
    .C(_01235_),
    .Y(_01236_));
 sky130_fd_sc_hd__a21o_1 _19401_ (.A1(_01234_),
    .A2(_01235_),
    .B1(_01229_),
    .X(_01237_));
 sky130_fd_sc_hd__a22o_1 _19402_ (.A1(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[4] ),
    .A2(net192),
    .B1(net247),
    .B2(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[3] ),
    .X(_01238_));
 sky130_fd_sc_hd__nand4_4 _19403_ (.A(_11697_),
    .B(_11693_),
    .C(net190),
    .D(_11687_),
    .Y(_01239_));
 sky130_fd_sc_hd__nand4_4 _19404_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[2] ),
    .B(_11692_),
    .C(_01238_),
    .D(_01239_),
    .Y(_01240_));
 sky130_fd_sc_hd__a22o_1 _19405_ (.A1(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[2] ),
    .A2(_11692_),
    .B1(_01238_),
    .B2(_01239_),
    .X(_01241_));
 sky130_fd_sc_hd__and4_1 _19406_ (.A(_11701_),
    .B(_11677_),
    .C(_01240_),
    .D(_01241_),
    .X(_01242_));
 sky130_fd_sc_hd__a22oi_1 _19407_ (.A1(_11701_),
    .A2(_11677_),
    .B1(_01240_),
    .B2(_01241_),
    .Y(_01243_));
 sky130_fd_sc_hd__nor2_1 _19408_ (.A(_01242_),
    .B(_01243_),
    .Y(_01244_));
 sky130_fd_sc_hd__and3_1 _19409_ (.A(_01236_),
    .B(_01237_),
    .C(_01244_),
    .X(_01245_));
 sky130_fd_sc_hd__a21oi_1 _19410_ (.A1(_01236_),
    .A2(_01237_),
    .B1(_01244_),
    .Y(_01246_));
 sky130_fd_sc_hd__nor3b_4 _19411_ (.A(_01245_),
    .B(_01246_),
    .C_N(_01218_),
    .Y(_01247_));
 sky130_fd_sc_hd__o21ba_1 _19412_ (.A1(_01245_),
    .A2(_01246_),
    .B1_N(_01218_),
    .X(_01248_));
 sky130_fd_sc_hd__nand2_1 _19413_ (.A(_01207_),
    .B(_01210_),
    .Y(_01249_));
 sky130_fd_sc_hd__or3b_4 _19414_ (.A(_01247_),
    .B(_01248_),
    .C_N(_01249_),
    .X(_01250_));
 sky130_fd_sc_hd__o21bai_2 _19415_ (.A1(_01247_),
    .A2(_01248_),
    .B1_N(_01249_),
    .Y(_01251_));
 sky130_fd_sc_hd__nor3b_1 _19416_ (.A(_01218_),
    .B(_01219_),
    .C_N(_01220_),
    .Y(_01252_));
 sky130_fd_sc_hd__a21o_1 _19417_ (.A1(_01195_),
    .A2(_01222_),
    .B1(_01252_),
    .X(_01253_));
 sky130_fd_sc_hd__nand3_1 _19418_ (.A(_01250_),
    .B(_01251_),
    .C(_01253_),
    .Y(_01254_));
 sky130_fd_sc_hd__a21o_1 _19419_ (.A1(_01250_),
    .A2(_01251_),
    .B1(_01253_),
    .X(_01255_));
 sky130_fd_sc_hd__and3_1 _19420_ (.A(_01228_),
    .B(_01254_),
    .C(_01255_),
    .X(_01256_));
 sky130_fd_sc_hd__a21o_1 _19421_ (.A1(_01254_),
    .A2(_01255_),
    .B1(_01228_),
    .X(_01257_));
 sky130_fd_sc_hd__and3b_1 _19422_ (.A_N(_01256_),
    .B(_01257_),
    .C(_06168_),
    .X(_01258_));
 sky130_fd_sc_hd__o21a_1 _19423_ (.A1(_01227_),
    .A2(_01258_),
    .B1(_04870_),
    .X(_00731_));
 sky130_fd_sc_hd__nand2_1 _19424_ (.A(_01250_),
    .B(_01251_),
    .Y(_01259_));
 sky130_fd_sc_hd__nor3b_1 _19425_ (.A(_01247_),
    .B(_01248_),
    .C_N(_01249_),
    .Y(_01260_));
 sky130_fd_sc_hd__a21bo_1 _19426_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[5] ),
    .A2(_01230_),
    .B1_N(_01231_),
    .X(_01261_));
 sky130_fd_sc_hd__a22o_1 _19427_ (.A1(_11683_),
    .A2(net195),
    .B1(_11704_),
    .B2(_11678_),
    .X(_01262_));
 sky130_fd_sc_hd__nand4_1 _19428_ (.A(_11683_),
    .B(_11678_),
    .C(_11700_),
    .D(_11705_),
    .Y(_01263_));
 sky130_fd_sc_hd__and3_1 _19429_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[6] ),
    .B(_01262_),
    .C(_01263_),
    .X(_01264_));
 sky130_fd_sc_hd__a21oi_2 _19430_ (.A1(net231),
    .A2(_01263_),
    .B1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[6] ),
    .Y(_01265_));
 sky130_fd_sc_hd__a211o_1 _19431_ (.A1(_01239_),
    .A2(_01240_),
    .B1(_01264_),
    .C1(_01265_),
    .X(_01266_));
 sky130_fd_sc_hd__o211ai_2 _19432_ (.A1(_01264_),
    .A2(_01265_),
    .B1(_01239_),
    .C1(_01240_),
    .Y(_01267_));
 sky130_fd_sc_hd__nand3_2 _19433_ (.A(_01261_),
    .B(net232),
    .C(_01267_),
    .Y(_01268_));
 sky130_fd_sc_hd__a21o_1 _19434_ (.A1(_01266_),
    .A2(_01267_),
    .B1(_01261_),
    .X(_01269_));
 sky130_fd_sc_hd__a22o_1 _19435_ (.A1(_11697_),
    .A2(_11687_),
    .B1(_11692_),
    .B2(_11693_),
    .X(_01270_));
 sky130_fd_sc_hd__nand4_2 _19436_ (.A(_11697_),
    .B(_11693_),
    .C(_11687_),
    .D(_11692_),
    .Y(_01271_));
 sky130_fd_sc_hd__nand4_2 _19437_ (.A(_11688_),
    .B(_11696_),
    .C(_01270_),
    .D(_01271_),
    .Y(_01272_));
 sky130_fd_sc_hd__a22o_1 _19438_ (.A1(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[2] ),
    .A2(_11696_),
    .B1(_01270_),
    .B2(_01271_),
    .X(_01273_));
 sky130_fd_sc_hd__a22oi_1 _19439_ (.A1(_11703_),
    .A2(net244),
    .B1(_11682_),
    .B2(_11701_),
    .Y(_01274_));
 sky130_fd_sc_hd__and4_1 _19440_ (.A(_11703_),
    .B(_11701_),
    .C(net243),
    .D(_11682_),
    .X(_01275_));
 sky130_fd_sc_hd__nor2_1 _19441_ (.A(_01274_),
    .B(_01275_),
    .Y(_01276_));
 sky130_fd_sc_hd__nand3_1 _19442_ (.A(_01272_),
    .B(_01273_),
    .C(_01276_),
    .Y(_01277_));
 sky130_fd_sc_hd__a21o_1 _19443_ (.A1(_01272_),
    .A2(_01273_),
    .B1(_01276_),
    .X(_01278_));
 sky130_fd_sc_hd__nand3_1 _19444_ (.A(_01242_),
    .B(_01277_),
    .C(_01278_),
    .Y(_01279_));
 sky130_fd_sc_hd__a21o_1 _19445_ (.A1(_01277_),
    .A2(_01278_),
    .B1(_01242_),
    .X(_01280_));
 sky130_fd_sc_hd__nand4_2 _19446_ (.A(_01268_),
    .B(_01269_),
    .C(_01279_),
    .D(_01280_),
    .Y(_01281_));
 sky130_fd_sc_hd__a22o_1 _19447_ (.A1(_01268_),
    .A2(_01269_),
    .B1(_01279_),
    .B2(_01280_),
    .X(_01282_));
 sky130_fd_sc_hd__and3_1 _19448_ (.A(_01245_),
    .B(_01281_),
    .C(_01282_),
    .X(_01283_));
 sky130_fd_sc_hd__a21oi_1 _19449_ (.A1(_01281_),
    .A2(net236),
    .B1(_01245_),
    .Y(_01284_));
 sky130_fd_sc_hd__a211o_1 _19450_ (.A1(net218),
    .A2(_01236_),
    .B1(_01283_),
    .C1(_01284_),
    .X(_01285_));
 sky130_fd_sc_hd__o211ai_2 _19451_ (.A1(_01283_),
    .A2(_01284_),
    .B1(net218),
    .C1(_01236_),
    .Y(_01286_));
 sky130_fd_sc_hd__o211a_1 _19452_ (.A1(_01247_),
    .A2(_01260_),
    .B1(_01285_),
    .C1(_01286_),
    .X(_01287_));
 sky130_fd_sc_hd__a211oi_1 _19453_ (.A1(net237),
    .A2(_01286_),
    .B1(_01247_),
    .C1(_01260_),
    .Y(_01288_));
 sky130_fd_sc_hd__or4_1 _19454_ (.A(_01221_),
    .B(_01259_),
    .C(_01287_),
    .D(_01288_),
    .X(_01289_));
 sky130_fd_sc_hd__o22ai_2 _19455_ (.A1(_01221_),
    .A2(_01259_),
    .B1(_01287_),
    .B2(_01288_),
    .Y(_01290_));
 sky130_fd_sc_hd__nand2_1 _19456_ (.A(_01289_),
    .B(_01290_),
    .Y(_01291_));
 sky130_fd_sc_hd__and3_1 _19457_ (.A(_01195_),
    .B(_01221_),
    .C(_01222_),
    .X(_01292_));
 sky130_fd_sc_hd__a31o_1 _19458_ (.A1(_01250_),
    .A2(_01251_),
    .A3(_01292_),
    .B1(_01256_),
    .X(_01293_));
 sky130_fd_sc_hd__xnor2_2 _19459_ (.A(_01291_),
    .B(_01293_),
    .Y(_01294_));
 sky130_fd_sc_hd__mux2_1 _19460_ (.A0(\top_inst.deskew_buff_inst.col_input[6] ),
    .A1(_01294_),
    .S(_08307_),
    .X(_01295_));
 sky130_fd_sc_hd__and2_1 _19461_ (.A(_11722_),
    .B(_01295_),
    .X(_01296_));
 sky130_fd_sc_hd__clkbuf_1 _19462_ (.A(_01296_),
    .X(_00732_));
 sky130_fd_sc_hd__inv_2 _19463_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[7] ),
    .Y(_01297_));
 sky130_fd_sc_hd__buf_2 _19464_ (.A(_01297_),
    .X(_01298_));
 sky130_fd_sc_hd__a21boi_1 _19465_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[6] ),
    .A2(net231),
    .B1_N(_01263_),
    .Y(_01299_));
 sky130_fd_sc_hd__nand2_1 _19466_ (.A(_01271_),
    .B(_01272_),
    .Y(_01300_));
 sky130_fd_sc_hd__and3_1 _19467_ (.A(_11678_),
    .B(_11705_),
    .C(_11708_),
    .X(_01301_));
 sky130_fd_sc_hd__a22o_1 _19468_ (.A1(_11683_),
    .A2(_11704_),
    .B1(_11708_),
    .B2(_11678_),
    .X(_01302_));
 sky130_fd_sc_hd__a21bo_1 _19469_ (.A1(_11684_),
    .A2(_01301_),
    .B1_N(_01302_),
    .X(_01303_));
 sky130_fd_sc_hd__xor2_2 _19470_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[7] ),
    .B(_01303_),
    .X(_01304_));
 sky130_fd_sc_hd__xnor2_1 _19471_ (.A(_01300_),
    .B(_01304_),
    .Y(_01305_));
 sky130_fd_sc_hd__xnor2_1 _19472_ (.A(_01299_),
    .B(_01305_),
    .Y(_01306_));
 sky130_fd_sc_hd__and3_1 _19473_ (.A(_01272_),
    .B(_01273_),
    .C(_01276_),
    .X(_01307_));
 sky130_fd_sc_hd__nand2_1 _19474_ (.A(_11688_),
    .B(_11700_),
    .Y(_01308_));
 sky130_fd_sc_hd__a22oi_1 _19475_ (.A1(_11697_),
    .A2(_11692_),
    .B1(_11696_),
    .B2(_11693_),
    .Y(_01309_));
 sky130_fd_sc_hd__and4_1 _19476_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[3] ),
    .C(net239),
    .D(_11696_),
    .X(_01310_));
 sky130_fd_sc_hd__nor2_1 _19477_ (.A(_01309_),
    .B(_01310_),
    .Y(_01311_));
 sky130_fd_sc_hd__xnor2_1 _19478_ (.A(_01308_),
    .B(_01311_),
    .Y(_01312_));
 sky130_fd_sc_hd__and2_1 _19479_ (.A(_11701_),
    .B(net248),
    .X(_01313_));
 sky130_fd_sc_hd__inv_2 _19480_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[6] ),
    .Y(_01314_));
 sky130_fd_sc_hd__or4b_4 _19481_ (.A(_01297_),
    .B(_01314_),
    .C(_11676_),
    .D_N(net189),
    .X(_01315_));
 sky130_fd_sc_hd__a2bb2o_1 _19482_ (.A1_N(_01298_),
    .A2_N(net242),
    .B1(net190),
    .B2(_11703_),
    .X(_01316_));
 sky130_fd_sc_hd__nand3_1 _19483_ (.A(_01313_),
    .B(_01315_),
    .C(_01316_),
    .Y(_01317_));
 sky130_fd_sc_hd__a21o_1 _19484_ (.A1(_01315_),
    .A2(_01316_),
    .B1(_01313_),
    .X(_01318_));
 sky130_fd_sc_hd__nand3_1 _19485_ (.A(_01275_),
    .B(_01317_),
    .C(_01318_),
    .Y(_01319_));
 sky130_fd_sc_hd__a21o_1 _19486_ (.A1(_01317_),
    .A2(_01318_),
    .B1(_01275_),
    .X(_01320_));
 sky130_fd_sc_hd__nand3_1 _19487_ (.A(_01312_),
    .B(_01319_),
    .C(_01320_),
    .Y(_01321_));
 sky130_fd_sc_hd__a21o_1 _19488_ (.A1(_01319_),
    .A2(_01320_),
    .B1(_01312_),
    .X(_01322_));
 sky130_fd_sc_hd__nand3_2 _19489_ (.A(_01307_),
    .B(_01321_),
    .C(_01322_),
    .Y(_01323_));
 sky130_fd_sc_hd__a21o_1 _19490_ (.A1(_01321_),
    .A2(_01322_),
    .B1(_01307_),
    .X(_01324_));
 sky130_fd_sc_hd__nand3_1 _19491_ (.A(_01306_),
    .B(_01323_),
    .C(_01324_),
    .Y(_01325_));
 sky130_fd_sc_hd__a21o_1 _19492_ (.A1(_01323_),
    .A2(_01324_),
    .B1(_01306_),
    .X(_01326_));
 sky130_fd_sc_hd__nand2_1 _19493_ (.A(_01279_),
    .B(_01281_),
    .Y(_01327_));
 sky130_fd_sc_hd__and3_1 _19494_ (.A(_01325_),
    .B(_01326_),
    .C(_01327_),
    .X(_01328_));
 sky130_fd_sc_hd__a21oi_1 _19495_ (.A1(_01325_),
    .A2(_01326_),
    .B1(_01327_),
    .Y(_01329_));
 sky130_fd_sc_hd__a211oi_2 _19496_ (.A1(net197),
    .A2(_01268_),
    .B1(_01328_),
    .C1(_01329_),
    .Y(_01330_));
 sky130_fd_sc_hd__o211a_1 _19497_ (.A1(_01328_),
    .A2(_01329_),
    .B1(net198),
    .C1(_01268_),
    .X(_01331_));
 sky130_fd_sc_hd__and2b_1 _19498_ (.A_N(_01283_),
    .B(_01285_),
    .X(_01332_));
 sky130_fd_sc_hd__nor3_2 _19499_ (.A(net241),
    .B(_01331_),
    .C(_01332_),
    .Y(_01333_));
 sky130_fd_sc_hd__o21ai_2 _19500_ (.A1(_01330_),
    .A2(_01331_),
    .B1(_01332_),
    .Y(_01334_));
 sky130_fd_sc_hd__or3b_1 _19501_ (.A(_01298_),
    .B(_01333_),
    .C_N(_01334_),
    .X(_01335_));
 sky130_fd_sc_hd__or3_4 _19502_ (.A(net241),
    .B(_01331_),
    .C(_01332_),
    .X(_01336_));
 sky130_fd_sc_hd__a21o_1 _19503_ (.A1(_01336_),
    .A2(_01334_),
    .B1(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[7] ),
    .X(_01337_));
 sky130_fd_sc_hd__and3_1 _19504_ (.A(_01287_),
    .B(_01335_),
    .C(_01337_),
    .X(_01338_));
 sky130_fd_sc_hd__a21o_1 _19505_ (.A1(_01335_),
    .A2(_01337_),
    .B1(_01287_),
    .X(_01339_));
 sky130_fd_sc_hd__or2b_1 _19506_ (.A(_01338_),
    .B_N(_01339_),
    .X(_01340_));
 sky130_fd_sc_hd__a21bo_2 _19507_ (.A1(_01290_),
    .A2(_01293_),
    .B1_N(_01289_),
    .X(_01341_));
 sky130_fd_sc_hd__xnor2_2 _19508_ (.A(_01340_),
    .B(_01341_),
    .Y(_01342_));
 sky130_fd_sc_hd__mux2_1 _19509_ (.A0(\top_inst.deskew_buff_inst.col_input[7] ),
    .A1(_01342_),
    .S(_08307_),
    .X(_01343_));
 sky130_fd_sc_hd__and2_1 _19510_ (.A(_11722_),
    .B(_01343_),
    .X(_01344_));
 sky130_fd_sc_hd__clkbuf_1 _19511_ (.A(_01344_),
    .X(_00733_));
 sky130_fd_sc_hd__a21oi_4 _19512_ (.A1(_01339_),
    .A2(_01341_),
    .B1(_01338_),
    .Y(_01345_));
 sky130_fd_sc_hd__nor2_1 _19513_ (.A(_01328_),
    .B(_01330_),
    .Y(_01346_));
 sky130_fd_sc_hd__or2b_1 _19514_ (.A(_01304_),
    .B_N(_01300_),
    .X(_01347_));
 sky130_fd_sc_hd__or2b_1 _19515_ (.A(_01299_),
    .B_N(_01305_),
    .X(_01348_));
 sky130_fd_sc_hd__nand2_1 _19516_ (.A(_01347_),
    .B(_01348_),
    .Y(_01349_));
 sky130_fd_sc_hd__a22o_1 _19517_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[7] ),
    .A2(_01302_),
    .B1(_01301_),
    .B2(_11684_),
    .X(_01350_));
 sky130_fd_sc_hd__a31o_1 _19518_ (.A1(_11688_),
    .A2(_11700_),
    .A3(_01311_),
    .B1(_01310_),
    .X(_01351_));
 sky130_fd_sc_hd__o21ai_4 _19519_ (.A1(_11683_),
    .A2(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[0] ),
    .B1(_11708_),
    .Y(_01352_));
 sky130_fd_sc_hd__and3_2 _19520_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[1] ),
    .B(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[0] ),
    .C(_11707_),
    .X(_01353_));
 sky130_fd_sc_hd__nor2_2 _19521_ (.A(_01352_),
    .B(_01353_),
    .Y(_01354_));
 sky130_fd_sc_hd__xnor2_1 _19522_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[8] ),
    .B(_01354_),
    .Y(_01355_));
 sky130_fd_sc_hd__xnor2_1 _19523_ (.A(_01351_),
    .B(_01355_),
    .Y(_01356_));
 sky130_fd_sc_hd__xor2_1 _19524_ (.A(_01350_),
    .B(_01356_),
    .X(_01357_));
 sky130_fd_sc_hd__nand2_1 _19525_ (.A(_11688_),
    .B(_11705_),
    .Y(_01358_));
 sky130_fd_sc_hd__a22oi_1 _19526_ (.A1(_11697_),
    .A2(_11696_),
    .B1(_11700_),
    .B2(_11693_),
    .Y(_01359_));
 sky130_fd_sc_hd__and4_1 _19527_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[3] ),
    .C(_11695_),
    .D(net195),
    .X(_01360_));
 sky130_fd_sc_hd__nor2_1 _19528_ (.A(_01359_),
    .B(_01360_),
    .Y(_01361_));
 sky130_fd_sc_hd__xnor2_2 _19529_ (.A(_01358_),
    .B(_01361_),
    .Y(_01362_));
 sky130_fd_sc_hd__and2_1 _19530_ (.A(_11701_),
    .B(_11692_),
    .X(_01363_));
 sky130_fd_sc_hd__or4b_4 _19531_ (.A(_01297_),
    .B(_01314_),
    .C(_11681_),
    .D_N(net246),
    .X(_01364_));
 sky130_fd_sc_hd__a2bb2o_2 _19532_ (.A1_N(_01298_),
    .A2_N(net190),
    .B1(net247),
    .B2(_11703_),
    .X(_01365_));
 sky130_fd_sc_hd__nand3_1 _19533_ (.A(_01363_),
    .B(_01364_),
    .C(_01365_),
    .Y(_01366_));
 sky130_fd_sc_hd__a21o_1 _19534_ (.A1(_01364_),
    .A2(_01365_),
    .B1(_01363_),
    .X(_01367_));
 sky130_fd_sc_hd__a21bo_1 _19535_ (.A1(_01313_),
    .A2(_01316_),
    .B1_N(_01315_),
    .X(_01368_));
 sky130_fd_sc_hd__nand3_1 _19536_ (.A(_01366_),
    .B(_01367_),
    .C(_01368_),
    .Y(_01369_));
 sky130_fd_sc_hd__a21o_1 _19537_ (.A1(_01366_),
    .A2(_01367_),
    .B1(_01368_),
    .X(_01370_));
 sky130_fd_sc_hd__nand3_1 _19538_ (.A(_01362_),
    .B(_01369_),
    .C(_01370_),
    .Y(_01371_));
 sky130_fd_sc_hd__a21o_1 _19539_ (.A1(_01369_),
    .A2(_01370_),
    .B1(_01362_),
    .X(_01372_));
 sky130_fd_sc_hd__a21bo_1 _19540_ (.A1(_01312_),
    .A2(_01320_),
    .B1_N(_01319_),
    .X(_01373_));
 sky130_fd_sc_hd__nand3_2 _19541_ (.A(_01371_),
    .B(_01372_),
    .C(_01373_),
    .Y(_01374_));
 sky130_fd_sc_hd__a21o_1 _19542_ (.A1(_01371_),
    .A2(_01372_),
    .B1(_01373_),
    .X(_01375_));
 sky130_fd_sc_hd__and3_1 _19543_ (.A(_01357_),
    .B(_01374_),
    .C(_01375_),
    .X(_01376_));
 sky130_fd_sc_hd__a21oi_1 _19544_ (.A1(_01374_),
    .A2(_01375_),
    .B1(_01357_),
    .Y(_01377_));
 sky130_fd_sc_hd__a211oi_2 _19545_ (.A1(_01323_),
    .A2(_01325_),
    .B1(_01376_),
    .C1(_01377_),
    .Y(_01378_));
 sky130_fd_sc_hd__o211a_1 _19546_ (.A1(_01376_),
    .A2(_01377_),
    .B1(_01323_),
    .C1(_01325_),
    .X(_01379_));
 sky130_fd_sc_hd__nor2_2 _19547_ (.A(_01378_),
    .B(_01379_),
    .Y(_01380_));
 sky130_fd_sc_hd__xor2_2 _19548_ (.A(_01349_),
    .B(_01380_),
    .X(_01381_));
 sky130_fd_sc_hd__xnor2_2 _19549_ (.A(_01346_),
    .B(_01381_),
    .Y(_01382_));
 sky130_fd_sc_hd__a21o_1 _19550_ (.A1(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[7] ),
    .A2(_01334_),
    .B1(_01333_),
    .X(_01383_));
 sky130_fd_sc_hd__xnor2_2 _19551_ (.A(_01382_),
    .B(_01383_),
    .Y(_01384_));
 sky130_fd_sc_hd__xor2_2 _19552_ (.A(_01345_),
    .B(net210),
    .X(_01385_));
 sky130_fd_sc_hd__clkbuf_4 _19553_ (.A(_06701_),
    .X(_01386_));
 sky130_fd_sc_hd__or2_1 _19554_ (.A(net846),
    .B(_01386_),
    .X(_01387_));
 sky130_fd_sc_hd__o211a_1 _19555_ (.A1(_11177_),
    .A2(_01385_),
    .B1(_01387_),
    .C1(_11714_),
    .X(_00734_));
 sky130_fd_sc_hd__nand2_1 _19556_ (.A(_01382_),
    .B(_01383_),
    .Y(_01388_));
 sky130_fd_sc_hd__o21ai_2 _19557_ (.A1(_01345_),
    .A2(_01384_),
    .B1(_01388_),
    .Y(_01389_));
 sky130_fd_sc_hd__or2b_4 _19558_ (.A(_01346_),
    .B_N(_01381_),
    .X(_01390_));
 sky130_fd_sc_hd__and2b_1 _19559_ (.A_N(_01355_),
    .B(_01351_),
    .X(_01391_));
 sky130_fd_sc_hd__a21o_1 _19560_ (.A1(_01350_),
    .A2(_01356_),
    .B1(_01391_),
    .X(_01392_));
 sky130_fd_sc_hd__nand3_1 _19561_ (.A(_01357_),
    .B(_01374_),
    .C(_01375_),
    .Y(_01393_));
 sky130_fd_sc_hd__o21a_1 _19562_ (.A1(_11684_),
    .A2(_11679_),
    .B1(_11709_),
    .X(_01394_));
 sky130_fd_sc_hd__buf_2 _19563_ (.A(_01394_),
    .X(_01395_));
 sky130_fd_sc_hd__clkbuf_4 _19564_ (.A(_01353_),
    .X(_01396_));
 sky130_fd_sc_hd__a21o_1 _19565_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[8] ),
    .A2(_01395_),
    .B1(_01396_),
    .X(_01397_));
 sky130_fd_sc_hd__a31o_1 _19566_ (.A1(_11688_),
    .A2(_11705_),
    .A3(_01361_),
    .B1(_01360_),
    .X(_01398_));
 sky130_fd_sc_hd__xnor2_2 _19567_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[9] ),
    .B(_01354_),
    .Y(_01399_));
 sky130_fd_sc_hd__xnor2_1 _19568_ (.A(_01398_),
    .B(_01399_),
    .Y(_01400_));
 sky130_fd_sc_hd__xor2_1 _19569_ (.A(_01397_),
    .B(_01400_),
    .X(_01401_));
 sky130_fd_sc_hd__nand2_4 _19570_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[2] ),
    .B(_11708_),
    .Y(_01402_));
 sky130_fd_sc_hd__and3_1 _19571_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[3] ),
    .C(_11700_),
    .X(_01403_));
 sky130_fd_sc_hd__a22o_1 _19572_ (.A1(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[4] ),
    .A2(net195),
    .B1(_11704_),
    .B2(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[3] ),
    .X(_01404_));
 sky130_fd_sc_hd__a21bo_1 _19573_ (.A1(_11705_),
    .A2(_01403_),
    .B1_N(_01404_),
    .X(_01405_));
 sky130_fd_sc_hd__xor2_2 _19574_ (.A(_01402_),
    .B(_01405_),
    .X(_01406_));
 sky130_fd_sc_hd__and2_1 _19575_ (.A(_11701_),
    .B(_11696_),
    .X(_01407_));
 sky130_fd_sc_hd__or4b_4 _19576_ (.A(_01297_),
    .B(_01314_),
    .C(_11686_),
    .D_N(net239),
    .X(_01408_));
 sky130_fd_sc_hd__a2bb2o_1 _19577_ (.A1_N(_01298_),
    .A2_N(_11686_),
    .B1(net239),
    .B2(_11703_),
    .X(_01409_));
 sky130_fd_sc_hd__nand3_1 _19578_ (.A(_01407_),
    .B(_01408_),
    .C(_01409_),
    .Y(_01410_));
 sky130_fd_sc_hd__a21o_1 _19579_ (.A1(_01408_),
    .A2(_01409_),
    .B1(_01407_),
    .X(_01411_));
 sky130_fd_sc_hd__a21bo_1 _19580_ (.A1(_01363_),
    .A2(_01365_),
    .B1_N(_01364_),
    .X(_01412_));
 sky130_fd_sc_hd__nand3_1 _19581_ (.A(_01410_),
    .B(_01411_),
    .C(_01412_),
    .Y(_01413_));
 sky130_fd_sc_hd__a21o_1 _19582_ (.A1(_01410_),
    .A2(_01411_),
    .B1(_01412_),
    .X(_01414_));
 sky130_fd_sc_hd__nand3_2 _19583_ (.A(_01406_),
    .B(_01413_),
    .C(_01414_),
    .Y(_01415_));
 sky130_fd_sc_hd__a21o_1 _19584_ (.A1(_01413_),
    .A2(_01414_),
    .B1(_01406_),
    .X(_01416_));
 sky130_fd_sc_hd__a21bo_1 _19585_ (.A1(_01362_),
    .A2(_01370_),
    .B1_N(_01369_),
    .X(_01417_));
 sky130_fd_sc_hd__nand3_4 _19586_ (.A(_01415_),
    .B(net1126),
    .C(_01417_),
    .Y(_01418_));
 sky130_fd_sc_hd__a21o_1 _19587_ (.A1(_01415_),
    .A2(_01416_),
    .B1(_01417_),
    .X(_01419_));
 sky130_fd_sc_hd__and3_1 _19588_ (.A(net249),
    .B(_01418_),
    .C(_01419_),
    .X(_01420_));
 sky130_fd_sc_hd__a21oi_1 _19589_ (.A1(_01418_),
    .A2(_01419_),
    .B1(net249),
    .Y(_01421_));
 sky130_fd_sc_hd__a211o_1 _19590_ (.A1(_01374_),
    .A2(_01393_),
    .B1(_01420_),
    .C1(_01421_),
    .X(_01422_));
 sky130_fd_sc_hd__o211ai_1 _19591_ (.A1(_01420_),
    .A2(_01421_),
    .B1(_01374_),
    .C1(_01393_),
    .Y(_01423_));
 sky130_fd_sc_hd__nand3_1 _19592_ (.A(_01392_),
    .B(_01422_),
    .C(_01423_),
    .Y(_01424_));
 sky130_fd_sc_hd__a21o_1 _19593_ (.A1(_01422_),
    .A2(_01423_),
    .B1(_01392_),
    .X(_01425_));
 sky130_fd_sc_hd__and2_1 _19594_ (.A(_01424_),
    .B(_01425_),
    .X(_01426_));
 sky130_fd_sc_hd__a21o_1 _19595_ (.A1(_01349_),
    .A2(_01380_),
    .B1(_01378_),
    .X(_01427_));
 sky130_fd_sc_hd__xnor2_2 _19596_ (.A(_01426_),
    .B(_01427_),
    .Y(_01428_));
 sky130_fd_sc_hd__xnor2_2 _19597_ (.A(_01390_),
    .B(_01428_),
    .Y(_01429_));
 sky130_fd_sc_hd__xnor2_2 _19598_ (.A(_01389_),
    .B(_01429_),
    .Y(_01430_));
 sky130_fd_sc_hd__or2_1 _19599_ (.A(net464),
    .B(_01386_),
    .X(_01431_));
 sky130_fd_sc_hd__o211a_1 _19600_ (.A1(_11177_),
    .A2(_01430_),
    .B1(_01431_),
    .C1(_11714_),
    .X(_00735_));
 sky130_fd_sc_hd__nand2_1 _19601_ (.A(_01426_),
    .B(_01427_),
    .Y(_01432_));
 sky130_fd_sc_hd__and2b_1 _19602_ (.A_N(_01399_),
    .B(_01398_),
    .X(_01433_));
 sky130_fd_sc_hd__a21o_1 _19603_ (.A1(_01397_),
    .A2(_01400_),
    .B1(_01433_),
    .X(_01434_));
 sky130_fd_sc_hd__nand3_1 _19604_ (.A(_01401_),
    .B(_01418_),
    .C(_01419_),
    .Y(_01435_));
 sky130_fd_sc_hd__a21o_1 _19605_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[9] ),
    .A2(_01395_),
    .B1(_01396_),
    .X(_01436_));
 sky130_fd_sc_hd__a32o_1 _19606_ (.A1(_11688_),
    .A2(_11709_),
    .A3(_01404_),
    .B1(_01403_),
    .B2(_11705_),
    .X(_01437_));
 sky130_fd_sc_hd__xnor2_1 _19607_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[10] ),
    .B(_01354_),
    .Y(_01438_));
 sky130_fd_sc_hd__xnor2_1 _19608_ (.A(_01437_),
    .B(_01438_),
    .Y(_01439_));
 sky130_fd_sc_hd__xor2_1 _19609_ (.A(_01436_),
    .B(_01439_),
    .X(_01440_));
 sky130_fd_sc_hd__and3_1 _19610_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[3] ),
    .B(_11704_),
    .C(_11708_),
    .X(_01441_));
 sky130_fd_sc_hd__a22o_1 _19611_ (.A1(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[4] ),
    .A2(_11704_),
    .B1(_11708_),
    .B2(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[3] ),
    .X(_01442_));
 sky130_fd_sc_hd__a21bo_1 _19612_ (.A1(_11697_),
    .A2(_01441_),
    .B1_N(_01442_),
    .X(_01443_));
 sky130_fd_sc_hd__xor2_1 _19613_ (.A(_01402_),
    .B(_01443_),
    .X(_01444_));
 sky130_fd_sc_hd__and2_1 _19614_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[5] ),
    .B(net195),
    .X(_01445_));
 sky130_fd_sc_hd__or4b_4 _19615_ (.A(_01297_),
    .B(_01314_),
    .C(_11691_),
    .D_N(_11695_),
    .X(_01446_));
 sky130_fd_sc_hd__a2bb2o_1 _19616_ (.A1_N(_01298_),
    .A2_N(_11691_),
    .B1(_11695_),
    .B2(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[6] ),
    .X(_01447_));
 sky130_fd_sc_hd__nand3_1 _19617_ (.A(_01445_),
    .B(_01446_),
    .C(_01447_),
    .Y(_01448_));
 sky130_fd_sc_hd__a21o_1 _19618_ (.A1(_01446_),
    .A2(_01447_),
    .B1(_01445_),
    .X(_01449_));
 sky130_fd_sc_hd__a21bo_1 _19619_ (.A1(_01407_),
    .A2(_01409_),
    .B1_N(_01408_),
    .X(_01450_));
 sky130_fd_sc_hd__nand3_1 _19620_ (.A(_01448_),
    .B(_01449_),
    .C(_01450_),
    .Y(_01451_));
 sky130_fd_sc_hd__a21o_1 _19621_ (.A1(_01448_),
    .A2(_01449_),
    .B1(_01450_),
    .X(_01452_));
 sky130_fd_sc_hd__nand3_1 _19622_ (.A(_01444_),
    .B(_01451_),
    .C(_01452_),
    .Y(_01453_));
 sky130_fd_sc_hd__a21o_1 _19623_ (.A1(_01451_),
    .A2(_01452_),
    .B1(_01444_),
    .X(_01454_));
 sky130_fd_sc_hd__a21bo_1 _19624_ (.A1(_01406_),
    .A2(_01414_),
    .B1_N(_01413_),
    .X(_01455_));
 sky130_fd_sc_hd__nand3_2 _19625_ (.A(_01453_),
    .B(_01454_),
    .C(_01455_),
    .Y(_01456_));
 sky130_fd_sc_hd__a21o_1 _19626_ (.A1(_01453_),
    .A2(_01454_),
    .B1(_01455_),
    .X(_01457_));
 sky130_fd_sc_hd__and3_1 _19627_ (.A(_01440_),
    .B(_01456_),
    .C(_01457_),
    .X(_01458_));
 sky130_fd_sc_hd__a21oi_1 _19628_ (.A1(_01456_),
    .A2(_01457_),
    .B1(_01440_),
    .Y(_01459_));
 sky130_fd_sc_hd__a211o_1 _19629_ (.A1(_01418_),
    .A2(_01435_),
    .B1(_01458_),
    .C1(_01459_),
    .X(_01460_));
 sky130_fd_sc_hd__o211ai_2 _19630_ (.A1(net196),
    .A2(_01459_),
    .B1(_01418_),
    .C1(_01435_),
    .Y(_01461_));
 sky130_fd_sc_hd__and3_1 _19631_ (.A(_01434_),
    .B(_01460_),
    .C(_01461_),
    .X(_01462_));
 sky130_fd_sc_hd__a21oi_1 _19632_ (.A1(_01460_),
    .A2(_01461_),
    .B1(_01434_),
    .Y(_01463_));
 sky130_fd_sc_hd__a211oi_2 _19633_ (.A1(_01422_),
    .A2(_01424_),
    .B1(net238),
    .C1(_01463_),
    .Y(_01464_));
 sky130_fd_sc_hd__o211a_1 _19634_ (.A1(_01462_),
    .A2(_01463_),
    .B1(_01422_),
    .C1(_01424_),
    .X(_01465_));
 sky130_fd_sc_hd__or2_4 _19635_ (.A(_01464_),
    .B(_01465_),
    .X(_01466_));
 sky130_fd_sc_hd__xnor2_1 _19636_ (.A(_01432_),
    .B(_01466_),
    .Y(_01467_));
 sky130_fd_sc_hd__a21boi_1 _19637_ (.A1(_01382_),
    .A2(_01383_),
    .B1_N(_01390_),
    .Y(_01468_));
 sky130_fd_sc_hd__o32a_1 _19638_ (.A1(_01345_),
    .A2(_01384_),
    .A3(_01429_),
    .B1(_01468_),
    .B2(_01428_),
    .X(_01469_));
 sky130_fd_sc_hd__or2_1 _19639_ (.A(_01467_),
    .B(_01469_),
    .X(_01470_));
 sky130_fd_sc_hd__a21oi_1 _19640_ (.A1(_01467_),
    .A2(_01469_),
    .B1(_05399_),
    .Y(_01471_));
 sky130_fd_sc_hd__a22o_1 _19641_ (.A1(\top_inst.deskew_buff_inst.col_input[10] ),
    .A2(_11723_),
    .B1(_01470_),
    .B2(_01471_),
    .X(_01472_));
 sky130_fd_sc_hd__and2_1 _19642_ (.A(_11722_),
    .B(_01472_),
    .X(_01473_));
 sky130_fd_sc_hd__clkbuf_1 _19643_ (.A(_01473_),
    .X(_00736_));
 sky130_fd_sc_hd__or2_1 _19644_ (.A(_01432_),
    .B(_01466_),
    .X(_01474_));
 sky130_fd_sc_hd__and2b_1 _19645_ (.A_N(_01438_),
    .B(_01437_),
    .X(_01475_));
 sky130_fd_sc_hd__a21o_1 _19646_ (.A1(_01436_),
    .A2(_01439_),
    .B1(_01475_),
    .X(_01476_));
 sky130_fd_sc_hd__nand3_1 _19647_ (.A(_01440_),
    .B(_01456_),
    .C(_01457_),
    .Y(_01477_));
 sky130_fd_sc_hd__a21o_1 _19648_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[10] ),
    .A2(_01395_),
    .B1(_01396_),
    .X(_01478_));
 sky130_fd_sc_hd__a32o_1 _19649_ (.A1(_11688_),
    .A2(_11709_),
    .A3(_01442_),
    .B1(_01441_),
    .B2(_11697_),
    .X(_01479_));
 sky130_fd_sc_hd__buf_4 _19650_ (.A(_01354_),
    .X(_01480_));
 sky130_fd_sc_hd__xnor2_1 _19651_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[11] ),
    .B(_01480_),
    .Y(_01481_));
 sky130_fd_sc_hd__xnor2_1 _19652_ (.A(_01479_),
    .B(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__xor2_1 _19653_ (.A(_01478_),
    .B(_01482_),
    .X(_01483_));
 sky130_fd_sc_hd__and3_1 _19654_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[3] ),
    .C(_11708_),
    .X(_01484_));
 sky130_fd_sc_hd__o21ai_2 _19655_ (.A1(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[4] ),
    .A2(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[3] ),
    .B1(_11709_),
    .Y(_01485_));
 sky130_fd_sc_hd__or3_4 _19656_ (.A(_01402_),
    .B(_01484_),
    .C(_01485_),
    .X(_01486_));
 sky130_fd_sc_hd__o21ai_4 _19657_ (.A1(_01484_),
    .A2(_01485_),
    .B1(_01402_),
    .Y(_01487_));
 sky130_fd_sc_hd__nand2_2 _19658_ (.A(_01486_),
    .B(_01487_),
    .Y(_01488_));
 sky130_fd_sc_hd__and2_1 _19659_ (.A(_11701_),
    .B(_11704_),
    .X(_01489_));
 sky130_fd_sc_hd__or4b_4 _19660_ (.A(_01297_),
    .B(_01314_),
    .C(_11695_),
    .D_N(net235),
    .X(_01490_));
 sky130_fd_sc_hd__a2bb2o_1 _19661_ (.A1_N(_01298_),
    .A2_N(_11695_),
    .B1(net194),
    .B2(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[6] ),
    .X(_01491_));
 sky130_fd_sc_hd__nand3_1 _19662_ (.A(_01489_),
    .B(_01490_),
    .C(_01491_),
    .Y(_01492_));
 sky130_fd_sc_hd__a21o_1 _19663_ (.A1(_01490_),
    .A2(_01491_),
    .B1(_01489_),
    .X(_01493_));
 sky130_fd_sc_hd__a21bo_1 _19664_ (.A1(_01445_),
    .A2(_01447_),
    .B1_N(_01446_),
    .X(_01494_));
 sky130_fd_sc_hd__and3_1 _19665_ (.A(_01492_),
    .B(_01493_),
    .C(_01494_),
    .X(_01495_));
 sky130_fd_sc_hd__a21oi_1 _19666_ (.A1(_01492_),
    .A2(_01493_),
    .B1(_01494_),
    .Y(_01496_));
 sky130_fd_sc_hd__or3_4 _19667_ (.A(_01488_),
    .B(_01495_),
    .C(_01496_),
    .X(_01497_));
 sky130_fd_sc_hd__o21ai_1 _19668_ (.A1(_01495_),
    .A2(_01496_),
    .B1(_01488_),
    .Y(_01498_));
 sky130_fd_sc_hd__a21bo_1 _19669_ (.A1(_01444_),
    .A2(_01452_),
    .B1_N(_01451_),
    .X(_01499_));
 sky130_fd_sc_hd__nand3_2 _19670_ (.A(_01497_),
    .B(_01498_),
    .C(_01499_),
    .Y(_01500_));
 sky130_fd_sc_hd__a21o_1 _19671_ (.A1(_01497_),
    .A2(_01498_),
    .B1(_01499_),
    .X(_01501_));
 sky130_fd_sc_hd__and3_1 _19672_ (.A(_01483_),
    .B(_01500_),
    .C(_01501_),
    .X(_01502_));
 sky130_fd_sc_hd__a21oi_1 _19673_ (.A1(_01500_),
    .A2(net250),
    .B1(_01483_),
    .Y(_01503_));
 sky130_fd_sc_hd__a211o_1 _19674_ (.A1(_01456_),
    .A2(_01477_),
    .B1(_01502_),
    .C1(_01503_),
    .X(_01504_));
 sky130_fd_sc_hd__o211ai_2 _19675_ (.A1(_01502_),
    .A2(_01503_),
    .B1(_01456_),
    .C1(_01477_),
    .Y(_01505_));
 sky130_fd_sc_hd__and3_1 _19676_ (.A(_01476_),
    .B(_01504_),
    .C(_01505_),
    .X(_01506_));
 sky130_fd_sc_hd__a21oi_1 _19677_ (.A1(_01504_),
    .A2(_01505_),
    .B1(_01476_),
    .Y(_01507_));
 sky130_fd_sc_hd__nor2_4 _19678_ (.A(_01506_),
    .B(_01507_),
    .Y(_01508_));
 sky130_fd_sc_hd__a21bo_1 _19679_ (.A1(_01434_),
    .A2(_01461_),
    .B1_N(_01460_),
    .X(_01509_));
 sky130_fd_sc_hd__xnor2_2 _19680_ (.A(_01508_),
    .B(_01509_),
    .Y(_01510_));
 sky130_fd_sc_hd__xnor2_2 _19681_ (.A(net1116),
    .B(_01510_),
    .Y(_01511_));
 sky130_fd_sc_hd__a21oi_1 _19682_ (.A1(_01474_),
    .A2(_01470_),
    .B1(_01511_),
    .Y(_01512_));
 sky130_fd_sc_hd__a31o_1 _19683_ (.A1(_01474_),
    .A2(_01470_),
    .A3(_01511_),
    .B1(_10957_),
    .X(_01513_));
 sky130_fd_sc_hd__o221a_1 _19684_ (.A1(net1092),
    .A2(_01202_),
    .B1(_01512_),
    .B2(_01513_),
    .C1(_11228_),
    .X(_00737_));
 sky130_fd_sc_hd__or4b_4 _19685_ (.A(_01384_),
    .B(_01429_),
    .C(_01467_),
    .D_N(_01511_),
    .X(_01514_));
 sky130_fd_sc_hd__or4b_4 _19686_ (.A(_01428_),
    .B(_01467_),
    .C(_01468_),
    .D_N(_01511_),
    .X(_01515_));
 sky130_fd_sc_hd__inv_2 _19687_ (.A(net253),
    .Y(_01516_));
 sky130_fd_sc_hd__a21o_1 _19688_ (.A1(_01516_),
    .A2(_01474_),
    .B1(_01510_),
    .X(_01517_));
 sky130_fd_sc_hd__o211a_4 _19689_ (.A1(_01345_),
    .A2(_01514_),
    .B1(_01515_),
    .C1(_01517_),
    .X(_01518_));
 sky130_fd_sc_hd__nand2_1 _19690_ (.A(_01508_),
    .B(_01509_),
    .Y(_01519_));
 sky130_fd_sc_hd__a21bo_1 _19691_ (.A1(_01476_),
    .A2(_01505_),
    .B1_N(_01504_),
    .X(_01520_));
 sky130_fd_sc_hd__and2b_1 _19692_ (.A_N(_01481_),
    .B(_01479_),
    .X(_01521_));
 sky130_fd_sc_hd__a21o_1 _19693_ (.A1(_01478_),
    .A2(_01482_),
    .B1(_01521_),
    .X(_01522_));
 sky130_fd_sc_hd__nand3_1 _19694_ (.A(_01483_),
    .B(_01500_),
    .C(net251),
    .Y(_01523_));
 sky130_fd_sc_hd__nand3_4 _19695_ (.A(_11684_),
    .B(_11679_),
    .C(_11709_),
    .Y(_01524_));
 sky130_fd_sc_hd__nand2_1 _19696_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[11] ),
    .B(_01480_),
    .Y(_01525_));
 sky130_fd_sc_hd__nand2_1 _19697_ (.A(_01524_),
    .B(_01525_),
    .Y(_01526_));
 sky130_fd_sc_hd__o21ba_1 _19698_ (.A1(_01402_),
    .A2(_01485_),
    .B1_N(_01484_),
    .X(_01527_));
 sky130_fd_sc_hd__buf_4 _19699_ (.A(_01527_),
    .X(_01528_));
 sky130_fd_sc_hd__xnor2_1 _19700_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[12] ),
    .B(_01480_),
    .Y(_01529_));
 sky130_fd_sc_hd__xor2_1 _19701_ (.A(_01528_),
    .B(_01529_),
    .X(_01530_));
 sky130_fd_sc_hd__xor2_1 _19702_ (.A(_01526_),
    .B(_01530_),
    .X(_01531_));
 sky130_fd_sc_hd__a21bo_1 _19703_ (.A1(_01489_),
    .A2(_01491_),
    .B1_N(_01490_),
    .X(_01532_));
 sky130_fd_sc_hd__and2_1 _19704_ (.A(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[5] ),
    .B(_11707_),
    .X(_01533_));
 sky130_fd_sc_hd__clkbuf_2 _19705_ (.A(_01533_),
    .X(_01534_));
 sky130_fd_sc_hd__or4b_4 _19706_ (.A(_01297_),
    .B(_01314_),
    .C(_11699_),
    .D_N(_11704_),
    .X(_01535_));
 sky130_fd_sc_hd__a2bb2o_1 _19707_ (.A1_N(_01298_),
    .A2_N(_11700_),
    .B1(_11705_),
    .B2(_11703_),
    .X(_01536_));
 sky130_fd_sc_hd__nand3_1 _19708_ (.A(_01534_),
    .B(_01535_),
    .C(_01536_),
    .Y(_01537_));
 sky130_fd_sc_hd__a21o_1 _19709_ (.A1(_01535_),
    .A2(_01536_),
    .B1(_01534_),
    .X(_01538_));
 sky130_fd_sc_hd__and3_1 _19710_ (.A(_01532_),
    .B(_01537_),
    .C(_01538_),
    .X(_01539_));
 sky130_fd_sc_hd__a21oi_1 _19711_ (.A1(_01537_),
    .A2(_01538_),
    .B1(_01532_),
    .Y(_01540_));
 sky130_fd_sc_hd__or3_1 _19712_ (.A(_01488_),
    .B(_01539_),
    .C(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__o21ai_1 _19713_ (.A1(_01539_),
    .A2(_01540_),
    .B1(_01488_),
    .Y(_01542_));
 sky130_fd_sc_hd__o21bai_1 _19714_ (.A1(_01488_),
    .A2(_01496_),
    .B1_N(_01495_),
    .Y(_01543_));
 sky130_fd_sc_hd__nand3_1 _19715_ (.A(_01541_),
    .B(_01542_),
    .C(_01543_),
    .Y(_01544_));
 sky130_fd_sc_hd__a21o_1 _19716_ (.A1(_01541_),
    .A2(_01542_),
    .B1(_01543_),
    .X(_01545_));
 sky130_fd_sc_hd__and3_1 _19717_ (.A(_01531_),
    .B(_01544_),
    .C(_01545_),
    .X(_01546_));
 sky130_fd_sc_hd__a21oi_1 _19718_ (.A1(_01544_),
    .A2(_01545_),
    .B1(_01531_),
    .Y(_01547_));
 sky130_fd_sc_hd__a211o_1 _19719_ (.A1(_01500_),
    .A2(_01523_),
    .B1(_01546_),
    .C1(_01547_),
    .X(_01548_));
 sky130_fd_sc_hd__o211ai_2 _19720_ (.A1(_01546_),
    .A2(_01547_),
    .B1(_01500_),
    .C1(_01523_),
    .Y(_01549_));
 sky130_fd_sc_hd__and3_1 _19721_ (.A(_01522_),
    .B(_01548_),
    .C(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__a21oi_1 _19722_ (.A1(_01548_),
    .A2(_01549_),
    .B1(_01522_),
    .Y(_01551_));
 sky130_fd_sc_hd__or2_1 _19723_ (.A(_01550_),
    .B(_01551_),
    .X(_01552_));
 sky130_fd_sc_hd__xor2_1 _19724_ (.A(_01520_),
    .B(_01552_),
    .X(_01553_));
 sky130_fd_sc_hd__or2_1 _19725_ (.A(_01519_),
    .B(_01553_),
    .X(_01554_));
 sky130_fd_sc_hd__nand2_1 _19726_ (.A(_01519_),
    .B(_01553_),
    .Y(_01555_));
 sky130_fd_sc_hd__nand2_2 _19727_ (.A(_01554_),
    .B(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__xor2_2 _19728_ (.A(_01518_),
    .B(_01556_),
    .X(_01557_));
 sky130_fd_sc_hd__or2_1 _19729_ (.A(net826),
    .B(_01386_),
    .X(_01558_));
 sky130_fd_sc_hd__o211a_1 _19730_ (.A1(_11177_),
    .A2(_01557_),
    .B1(_01558_),
    .C1(_11714_),
    .X(_00738_));
 sky130_fd_sc_hd__o21a_1 _19731_ (.A1(_01518_),
    .A2(_01556_),
    .B1(_01554_),
    .X(_01559_));
 sky130_fd_sc_hd__or2b_1 _19732_ (.A(_01552_),
    .B_N(_01520_),
    .X(_01560_));
 sky130_fd_sc_hd__clkbuf_4 _19733_ (.A(_01528_),
    .X(_01561_));
 sky130_fd_sc_hd__clkbuf_4 _19734_ (.A(_01561_),
    .X(_01562_));
 sky130_fd_sc_hd__clkbuf_4 _19735_ (.A(_01562_),
    .X(_01563_));
 sky130_fd_sc_hd__nor2_1 _19736_ (.A(_01563_),
    .B(_01529_),
    .Y(_01564_));
 sky130_fd_sc_hd__a21o_1 _19737_ (.A1(_01526_),
    .A2(_01530_),
    .B1(_01564_),
    .X(_01565_));
 sky130_fd_sc_hd__a21o_1 _19738_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[12] ),
    .A2(_01395_),
    .B1(_01396_),
    .X(_01566_));
 sky130_fd_sc_hd__xnor2_2 _19739_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[13] ),
    .B(_01480_),
    .Y(_01567_));
 sky130_fd_sc_hd__xor2_2 _19740_ (.A(_01528_),
    .B(_01567_),
    .X(_01568_));
 sky130_fd_sc_hd__xor2_2 _19741_ (.A(_01566_),
    .B(_01568_),
    .X(_01569_));
 sky130_fd_sc_hd__a21bo_1 _19742_ (.A1(_01534_),
    .A2(_01536_),
    .B1_N(_01535_),
    .X(_01570_));
 sky130_fd_sc_hd__or4b_1 _19743_ (.A(_01298_),
    .B(_01314_),
    .C(_11704_),
    .D_N(_11708_),
    .X(_01571_));
 sky130_fd_sc_hd__a2bb2o_1 _19744_ (.A1_N(_01298_),
    .A2_N(_11705_),
    .B1(_11708_),
    .B2(_11703_),
    .X(_01572_));
 sky130_fd_sc_hd__nand3_1 _19745_ (.A(_01534_),
    .B(_01571_),
    .C(_01572_),
    .Y(_01573_));
 sky130_fd_sc_hd__a21o_1 _19746_ (.A1(_01571_),
    .A2(_01572_),
    .B1(_01534_),
    .X(_01574_));
 sky130_fd_sc_hd__and3_1 _19747_ (.A(_01570_),
    .B(_01573_),
    .C(_01574_),
    .X(_01575_));
 sky130_fd_sc_hd__a21oi_1 _19748_ (.A1(_01573_),
    .A2(_01574_),
    .B1(_01570_),
    .Y(_01576_));
 sky130_fd_sc_hd__or3_1 _19749_ (.A(_01488_),
    .B(_01575_),
    .C(_01576_),
    .X(_01577_));
 sky130_fd_sc_hd__o21ai_1 _19750_ (.A1(_01575_),
    .A2(_01576_),
    .B1(_01488_),
    .Y(_01578_));
 sky130_fd_sc_hd__o21bai_1 _19751_ (.A1(_01488_),
    .A2(_01540_),
    .B1_N(_01539_),
    .Y(_01579_));
 sky130_fd_sc_hd__nand3_1 _19752_ (.A(_01577_),
    .B(_01578_),
    .C(_01579_),
    .Y(_01580_));
 sky130_fd_sc_hd__a21o_1 _19753_ (.A1(_01577_),
    .A2(_01578_),
    .B1(_01579_),
    .X(_01581_));
 sky130_fd_sc_hd__nand3_1 _19754_ (.A(_01569_),
    .B(_01580_),
    .C(_01581_),
    .Y(_01582_));
 sky130_fd_sc_hd__a21o_1 _19755_ (.A1(_01580_),
    .A2(_01581_),
    .B1(_01569_),
    .X(_01583_));
 sky130_fd_sc_hd__a21bo_1 _19756_ (.A1(_01531_),
    .A2(_01545_),
    .B1_N(_01544_),
    .X(_01584_));
 sky130_fd_sc_hd__and3_1 _19757_ (.A(_01582_),
    .B(_01583_),
    .C(_01584_),
    .X(_01585_));
 sky130_fd_sc_hd__a21oi_1 _19758_ (.A1(_01582_),
    .A2(_01583_),
    .B1(_01584_),
    .Y(_01586_));
 sky130_fd_sc_hd__nor2_2 _19759_ (.A(_01585_),
    .B(_01586_),
    .Y(_01587_));
 sky130_fd_sc_hd__xnor2_2 _19760_ (.A(_01565_),
    .B(_01587_),
    .Y(_01588_));
 sky130_fd_sc_hd__a21bo_1 _19761_ (.A1(_01522_),
    .A2(_01549_),
    .B1_N(_01548_),
    .X(_01589_));
 sky130_fd_sc_hd__xor2_2 _19762_ (.A(_01588_),
    .B(_01589_),
    .X(_01590_));
 sky130_fd_sc_hd__xnor2_2 _19763_ (.A(_01560_),
    .B(_01590_),
    .Y(_01591_));
 sky130_fd_sc_hd__xnor2_2 _19764_ (.A(_01559_),
    .B(_01591_),
    .Y(_01592_));
 sky130_fd_sc_hd__nand2_1 _19765_ (.A(_05317_),
    .B(_01592_),
    .Y(_01593_));
 sky130_fd_sc_hd__o211a_1 _19766_ (.A1(net596),
    .A2(_10616_),
    .B1(_01593_),
    .C1(_11714_),
    .X(_00739_));
 sky130_fd_sc_hd__a21oi_1 _19767_ (.A1(_01560_),
    .A2(_01554_),
    .B1(_01590_),
    .Y(_01594_));
 sky130_fd_sc_hd__nor3_1 _19768_ (.A(_01518_),
    .B(_01556_),
    .C(_01591_),
    .Y(_01595_));
 sky130_fd_sc_hd__or2b_1 _19769_ (.A(_01588_),
    .B_N(_01589_),
    .X(_01596_));
 sky130_fd_sc_hd__a21o_1 _19770_ (.A1(_01565_),
    .A2(_01587_),
    .B1(_01585_),
    .X(_01597_));
 sky130_fd_sc_hd__nor2_1 _19771_ (.A(_01562_),
    .B(_01567_),
    .Y(_01598_));
 sky130_fd_sc_hd__a21o_1 _19772_ (.A1(_01566_),
    .A2(_01568_),
    .B1(_01598_),
    .X(_01599_));
 sky130_fd_sc_hd__a21o_1 _19773_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[13] ),
    .A2(_01395_),
    .B1(_01396_),
    .X(_01600_));
 sky130_fd_sc_hd__xnor2_1 _19774_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[14] ),
    .B(_01480_),
    .Y(_01601_));
 sky130_fd_sc_hd__xor2_1 _19775_ (.A(_01528_),
    .B(_01601_),
    .X(_01602_));
 sky130_fd_sc_hd__xor2_1 _19776_ (.A(_01600_),
    .B(_01602_),
    .X(_01603_));
 sky130_fd_sc_hd__o21bai_2 _19777_ (.A1(_01488_),
    .A2(_01576_),
    .B1_N(_01575_),
    .Y(_01604_));
 sky130_fd_sc_hd__nor2_1 _19778_ (.A(_01298_),
    .B(_11709_),
    .Y(_01605_));
 sky130_fd_sc_hd__a211o_2 _19779_ (.A1(_11703_),
    .A2(_11709_),
    .B1(_01534_),
    .C1(_01605_),
    .X(_01606_));
 sky130_fd_sc_hd__a21boi_1 _19780_ (.A1(_01534_),
    .A2(_01572_),
    .B1_N(_01571_),
    .Y(_01607_));
 sky130_fd_sc_hd__and3_1 _19781_ (.A(_11703_),
    .B(_11701_),
    .C(_11709_),
    .X(_01608_));
 sky130_fd_sc_hd__o211a_1 _19782_ (.A1(_01607_),
    .A2(_01608_),
    .B1(_01486_),
    .C1(_01487_),
    .X(_01609_));
 sky130_fd_sc_hd__a211oi_2 _19783_ (.A1(_01486_),
    .A2(_01487_),
    .B1(_01607_),
    .C1(_01608_),
    .Y(_01610_));
 sky130_fd_sc_hd__a21oi_4 _19784_ (.A1(_01486_),
    .A2(_01487_),
    .B1(_01606_),
    .Y(_01611_));
 sky130_fd_sc_hd__a211o_1 _19785_ (.A1(_01606_),
    .A2(_01609_),
    .B1(_01610_),
    .C1(_01611_),
    .X(_01612_));
 sky130_fd_sc_hd__xnor2_1 _19786_ (.A(_01604_),
    .B(_01612_),
    .Y(_01613_));
 sky130_fd_sc_hd__xnor2_1 _19787_ (.A(_01603_),
    .B(_01613_),
    .Y(_01614_));
 sky130_fd_sc_hd__a21bo_1 _19788_ (.A1(_01569_),
    .A2(_01581_),
    .B1_N(_01580_),
    .X(_01615_));
 sky130_fd_sc_hd__xnor2_1 _19789_ (.A(_01614_),
    .B(_01615_),
    .Y(_01616_));
 sky130_fd_sc_hd__nand2_1 _19790_ (.A(_01599_),
    .B(_01616_),
    .Y(_01617_));
 sky130_fd_sc_hd__or2_1 _19791_ (.A(_01599_),
    .B(_01616_),
    .X(_01618_));
 sky130_fd_sc_hd__and2_1 _19792_ (.A(_01617_),
    .B(_01618_),
    .X(_01619_));
 sky130_fd_sc_hd__xnor2_1 _19793_ (.A(_01597_),
    .B(_01619_),
    .Y(_01620_));
 sky130_fd_sc_hd__xor2_1 _19794_ (.A(_01596_),
    .B(_01620_),
    .X(_01621_));
 sky130_fd_sc_hd__o21ai_1 _19795_ (.A1(_01594_),
    .A2(_01595_),
    .B1(_01621_),
    .Y(_01622_));
 sky130_fd_sc_hd__o31a_1 _19796_ (.A1(_01621_),
    .A2(_01594_),
    .A3(_01595_),
    .B1(_05311_),
    .X(_01623_));
 sky130_fd_sc_hd__a22o_1 _19797_ (.A1(\top_inst.deskew_buff_inst.col_input[14] ),
    .A2(_11723_),
    .B1(_01622_),
    .B2(_01623_),
    .X(_01624_));
 sky130_fd_sc_hd__and2_1 _19798_ (.A(_11722_),
    .B(_01624_),
    .X(_01625_));
 sky130_fd_sc_hd__clkbuf_1 _19799_ (.A(_01625_),
    .X(_00740_));
 sky130_fd_sc_hd__nor2_1 _19800_ (.A(_01596_),
    .B(_01620_),
    .Y(_01626_));
 sky130_fd_sc_hd__inv_2 _19801_ (.A(_01626_),
    .Y(_01627_));
 sky130_fd_sc_hd__and2_1 _19802_ (.A(_01597_),
    .B(_01619_),
    .X(_01628_));
 sky130_fd_sc_hd__or2b_1 _19803_ (.A(_01614_),
    .B_N(_01615_),
    .X(_01629_));
 sky130_fd_sc_hd__nor2_1 _19804_ (.A(_01562_),
    .B(_01601_),
    .Y(_01630_));
 sky130_fd_sc_hd__a21o_1 _19805_ (.A1(_01600_),
    .A2(_01602_),
    .B1(_01630_),
    .X(_01631_));
 sky130_fd_sc_hd__nor2_1 _19806_ (.A(_01611_),
    .B(_01610_),
    .Y(_01632_));
 sky130_fd_sc_hd__a21o_1 _19807_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[14] ),
    .A2(_01395_),
    .B1(_01396_),
    .X(_01633_));
 sky130_fd_sc_hd__xnor2_1 _19808_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[15] ),
    .B(_01480_),
    .Y(_01634_));
 sky130_fd_sc_hd__xor2_1 _19809_ (.A(_01528_),
    .B(_01634_),
    .X(_01635_));
 sky130_fd_sc_hd__xnor2_1 _19810_ (.A(_01633_),
    .B(_01635_),
    .Y(_01636_));
 sky130_fd_sc_hd__xnor2_1 _19811_ (.A(_01632_),
    .B(_01636_),
    .Y(_01637_));
 sky130_fd_sc_hd__nand2_1 _19812_ (.A(_01606_),
    .B(_01609_),
    .Y(_01638_));
 sky130_fd_sc_hd__a32o_1 _19813_ (.A1(_01604_),
    .A2(_01632_),
    .A3(_01638_),
    .B1(_01613_),
    .B2(_01603_),
    .X(_01639_));
 sky130_fd_sc_hd__xor2_1 _19814_ (.A(_01637_),
    .B(_01639_),
    .X(_01640_));
 sky130_fd_sc_hd__xnor2_1 _19815_ (.A(_01631_),
    .B(_01640_),
    .Y(_01641_));
 sky130_fd_sc_hd__a21oi_2 _19816_ (.A1(_01629_),
    .A2(_01617_),
    .B1(_01641_),
    .Y(_01642_));
 sky130_fd_sc_hd__and3_1 _19817_ (.A(_01629_),
    .B(_01617_),
    .C(_01641_),
    .X(_01643_));
 sky130_fd_sc_hd__nor2_1 _19818_ (.A(_01642_),
    .B(_01643_),
    .Y(_01644_));
 sky130_fd_sc_hd__xor2_1 _19819_ (.A(_01628_),
    .B(_01644_),
    .X(_01645_));
 sky130_fd_sc_hd__a21oi_1 _19820_ (.A1(_01627_),
    .A2(_01622_),
    .B1(_01645_),
    .Y(_01646_));
 sky130_fd_sc_hd__a31o_1 _19821_ (.A1(_01627_),
    .A2(_01622_),
    .A3(_01645_),
    .B1(_10957_),
    .X(_01647_));
 sky130_fd_sc_hd__o221a_1 _19822_ (.A1(net1093),
    .A2(_01202_),
    .B1(_01646_),
    .B2(_01647_),
    .C1(_11228_),
    .X(_00741_));
 sky130_fd_sc_hd__and2_1 _19823_ (.A(_01621_),
    .B(_01645_),
    .X(_01648_));
 sky130_fd_sc_hd__or3b_4 _19824_ (.A(_01556_),
    .B(_01591_),
    .C_N(_01648_),
    .X(_01649_));
 sky130_fd_sc_hd__o21a_1 _19825_ (.A1(_01628_),
    .A2(_01626_),
    .B1(_01644_),
    .X(_01650_));
 sky130_fd_sc_hd__a21oi_1 _19826_ (.A1(_01594_),
    .A2(_01648_),
    .B1(_01650_),
    .Y(_01651_));
 sky130_fd_sc_hd__o21ai_4 _19827_ (.A1(_01518_),
    .A2(_01649_),
    .B1(_01651_),
    .Y(_01652_));
 sky130_fd_sc_hd__and2_1 _19828_ (.A(_01637_),
    .B(_01639_),
    .X(_01653_));
 sky130_fd_sc_hd__a21o_1 _19829_ (.A1(_01631_),
    .A2(_01640_),
    .B1(_01653_),
    .X(_01654_));
 sky130_fd_sc_hd__nor2_1 _19830_ (.A(_01562_),
    .B(_01634_),
    .Y(_01655_));
 sky130_fd_sc_hd__a21o_1 _19831_ (.A1(_01633_),
    .A2(_01635_),
    .B1(_01655_),
    .X(_01656_));
 sky130_fd_sc_hd__o21ba_1 _19832_ (.A1(_01611_),
    .A2(_01636_),
    .B1_N(_01610_),
    .X(_01657_));
 sky130_fd_sc_hd__a21o_1 _19833_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[15] ),
    .A2(_01395_),
    .B1(_01396_),
    .X(_01658_));
 sky130_fd_sc_hd__or3b_1 _19834_ (.A(_01352_),
    .B(_01353_),
    .C_N(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[16] ),
    .X(_01659_));
 sky130_fd_sc_hd__a21o_1 _19835_ (.A1(_01394_),
    .A2(_01524_),
    .B1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[16] ),
    .X(_01660_));
 sky130_fd_sc_hd__nand3b_1 _19836_ (.A_N(_01528_),
    .B(_01659_),
    .C(_01660_),
    .Y(_01661_));
 sky130_fd_sc_hd__a21bo_1 _19837_ (.A1(_01659_),
    .A2(_01660_),
    .B1_N(_01528_),
    .X(_01662_));
 sky130_fd_sc_hd__nand3_1 _19838_ (.A(_01658_),
    .B(_01661_),
    .C(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__a21o_1 _19839_ (.A1(_01661_),
    .A2(_01662_),
    .B1(_01658_),
    .X(_01664_));
 sky130_fd_sc_hd__a21oi_1 _19840_ (.A1(_01663_),
    .A2(_01664_),
    .B1(_01611_),
    .Y(_01665_));
 sky130_fd_sc_hd__and3_1 _19841_ (.A(_01611_),
    .B(_01663_),
    .C(_01664_),
    .X(_01666_));
 sky130_fd_sc_hd__nor2_1 _19842_ (.A(_01665_),
    .B(_01666_),
    .Y(_01667_));
 sky130_fd_sc_hd__xnor2_1 _19843_ (.A(_01657_),
    .B(_01667_),
    .Y(_01668_));
 sky130_fd_sc_hd__xor2_1 _19844_ (.A(_01656_),
    .B(_01668_),
    .X(_01669_));
 sky130_fd_sc_hd__xnor2_1 _19845_ (.A(_01654_),
    .B(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__nand2_1 _19846_ (.A(_01642_),
    .B(_01670_),
    .Y(_01671_));
 sky130_fd_sc_hd__or2_1 _19847_ (.A(_01642_),
    .B(_01670_),
    .X(_01672_));
 sky130_fd_sc_hd__and2_1 _19848_ (.A(_01671_),
    .B(_01672_),
    .X(_01673_));
 sky130_fd_sc_hd__nand2_1 _19849_ (.A(_01652_),
    .B(_01673_),
    .Y(_01674_));
 sky130_fd_sc_hd__or2_1 _19850_ (.A(_01652_),
    .B(_01673_),
    .X(_01675_));
 sky130_fd_sc_hd__and2_1 _19851_ (.A(_01674_),
    .B(_01675_),
    .X(_01676_));
 sky130_fd_sc_hd__or2_1 _19852_ (.A(net311),
    .B(_01386_),
    .X(_01677_));
 sky130_fd_sc_hd__o211a_1 _19853_ (.A1(_11177_),
    .A2(_01676_),
    .B1(_01677_),
    .C1(_11714_),
    .X(_00742_));
 sky130_fd_sc_hd__or2b_1 _19854_ (.A(_01669_),
    .B_N(_01654_),
    .X(_01678_));
 sky130_fd_sc_hd__or2_1 _19855_ (.A(_01657_),
    .B(_01667_),
    .X(_01679_));
 sky130_fd_sc_hd__or2b_1 _19856_ (.A(_01668_),
    .B_N(_01656_),
    .X(_01680_));
 sky130_fd_sc_hd__nand2_1 _19857_ (.A(_01661_),
    .B(_01663_),
    .Y(_01681_));
 sky130_fd_sc_hd__and2_1 _19858_ (.A(_01524_),
    .B(_01659_),
    .X(_01682_));
 sky130_fd_sc_hd__or3b_1 _19859_ (.A(_01352_),
    .B(_01353_),
    .C_N(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[17] ),
    .X(_01683_));
 sky130_fd_sc_hd__a21o_1 _19860_ (.A1(_01394_),
    .A2(_01524_),
    .B1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[17] ),
    .X(_01684_));
 sky130_fd_sc_hd__nand3b_1 _19861_ (.A_N(_01527_),
    .B(_01683_),
    .C(_01684_),
    .Y(_01685_));
 sky130_fd_sc_hd__a21bo_1 _19862_ (.A1(_01683_),
    .A2(_01684_),
    .B1_N(_01527_),
    .X(_01686_));
 sky130_fd_sc_hd__nand2_1 _19863_ (.A(_01685_),
    .B(_01686_),
    .Y(_01687_));
 sky130_fd_sc_hd__xor2_2 _19864_ (.A(_01682_),
    .B(_01687_),
    .X(_01688_));
 sky130_fd_sc_hd__xnor2_1 _19865_ (.A(_01665_),
    .B(_01688_),
    .Y(_01689_));
 sky130_fd_sc_hd__xor2_1 _19866_ (.A(_01681_),
    .B(_01689_),
    .X(_01690_));
 sky130_fd_sc_hd__a21oi_2 _19867_ (.A1(_01679_),
    .A2(_01680_),
    .B1(_01690_),
    .Y(_01691_));
 sky130_fd_sc_hd__and3_1 _19868_ (.A(_01679_),
    .B(_01680_),
    .C(_01690_),
    .X(_01692_));
 sky130_fd_sc_hd__nor2_1 _19869_ (.A(_01691_),
    .B(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__xnor2_2 _19870_ (.A(_01678_),
    .B(_01693_),
    .Y(_01694_));
 sky130_fd_sc_hd__a21oi_1 _19871_ (.A1(_01671_),
    .A2(_01674_),
    .B1(_01694_),
    .Y(_01695_));
 sky130_fd_sc_hd__a31o_1 _19872_ (.A1(_01671_),
    .A2(_01674_),
    .A3(_01694_),
    .B1(_10957_),
    .X(_01696_));
 sky130_fd_sc_hd__o221a_1 _19873_ (.A1(net1096),
    .A2(_01202_),
    .B1(_01695_),
    .B2(_01696_),
    .C1(_11228_),
    .X(_00743_));
 sky130_fd_sc_hd__o21ai_2 _19874_ (.A1(_01682_),
    .A2(_01687_),
    .B1(_01685_),
    .Y(_01697_));
 sky130_fd_sc_hd__and2_1 _19875_ (.A(_01524_),
    .B(_01683_),
    .X(_01698_));
 sky130_fd_sc_hd__xnor2_2 _19876_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[18] ),
    .B(_01480_),
    .Y(_01699_));
 sky130_fd_sc_hd__xor2_2 _19877_ (.A(_01528_),
    .B(_01699_),
    .X(_01700_));
 sky130_fd_sc_hd__xnor2_2 _19878_ (.A(_01698_),
    .B(_01700_),
    .Y(_01701_));
 sky130_fd_sc_hd__or2_2 _19879_ (.A(_01611_),
    .B(_01688_),
    .X(_01702_));
 sky130_fd_sc_hd__xnor2_2 _19880_ (.A(_01701_),
    .B(_01702_),
    .Y(_01703_));
 sky130_fd_sc_hd__xnor2_2 _19881_ (.A(_01697_),
    .B(_01703_),
    .Y(_01704_));
 sky130_fd_sc_hd__nand2_1 _19882_ (.A(_01663_),
    .B(_01664_),
    .Y(_01705_));
 sky130_fd_sc_hd__or2b_1 _19883_ (.A(_01689_),
    .B_N(_01681_),
    .X(_01706_));
 sky130_fd_sc_hd__o21ai_2 _19884_ (.A1(_01705_),
    .A2(_01702_),
    .B1(_01706_),
    .Y(_01707_));
 sky130_fd_sc_hd__xnor2_2 _19885_ (.A(_01704_),
    .B(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hd__xor2_1 _19886_ (.A(_01691_),
    .B(_01708_),
    .X(_01709_));
 sky130_fd_sc_hd__a21boi_1 _19887_ (.A1(_01678_),
    .A2(_01671_),
    .B1_N(_01693_),
    .Y(_01710_));
 sky130_fd_sc_hd__a31oi_2 _19888_ (.A1(_01652_),
    .A2(_01673_),
    .A3(_01694_),
    .B1(_01710_),
    .Y(_01711_));
 sky130_fd_sc_hd__xnor2_1 _19889_ (.A(_01709_),
    .B(_01711_),
    .Y(_01712_));
 sky130_fd_sc_hd__mux2_1 _19890_ (.A0(\top_inst.deskew_buff_inst.col_input[18] ),
    .A1(_01712_),
    .S(_06140_),
    .X(_01713_));
 sky130_fd_sc_hd__and2_1 _19891_ (.A(_11722_),
    .B(_01713_),
    .X(_01714_));
 sky130_fd_sc_hd__clkbuf_1 _19892_ (.A(_01714_),
    .X(_00744_));
 sky130_fd_sc_hd__nor2_1 _19893_ (.A(_01691_),
    .B(_01708_),
    .Y(_01715_));
 sky130_fd_sc_hd__nand2_1 _19894_ (.A(_01691_),
    .B(_01708_),
    .Y(_01716_));
 sky130_fd_sc_hd__o21a_1 _19895_ (.A1(_01715_),
    .A2(_01711_),
    .B1(_01716_),
    .X(_01717_));
 sky130_fd_sc_hd__or2b_1 _19896_ (.A(_01704_),
    .B_N(_01707_),
    .X(_01718_));
 sky130_fd_sc_hd__or2b_1 _19897_ (.A(_01698_),
    .B_N(_01700_),
    .X(_01719_));
 sky130_fd_sc_hd__o21ai_2 _19898_ (.A1(_01562_),
    .A2(_01699_),
    .B1(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__a21o_2 _19899_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[18] ),
    .A2(_01395_),
    .B1(_01396_),
    .X(_01721_));
 sky130_fd_sc_hd__xnor2_1 _19900_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[19] ),
    .B(_01480_),
    .Y(_01722_));
 sky130_fd_sc_hd__nor2_1 _19901_ (.A(_01528_),
    .B(_01722_),
    .Y(_01723_));
 sky130_fd_sc_hd__nand2_1 _19902_ (.A(_01528_),
    .B(_01722_),
    .Y(_01724_));
 sky130_fd_sc_hd__and2b_1 _19903_ (.A_N(_01723_),
    .B(_01724_),
    .X(_01725_));
 sky130_fd_sc_hd__xor2_4 _19904_ (.A(_01721_),
    .B(_01725_),
    .X(_01726_));
 sky130_fd_sc_hd__nor2_1 _19905_ (.A(_01611_),
    .B(_01701_),
    .Y(_01727_));
 sky130_fd_sc_hd__xor2_2 _19906_ (.A(_01726_),
    .B(_01727_),
    .X(_01728_));
 sky130_fd_sc_hd__xnor2_2 _19907_ (.A(_01720_),
    .B(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__a22o_1 _19908_ (.A1(_01697_),
    .A2(_01703_),
    .B1(_01727_),
    .B2(_01688_),
    .X(_01730_));
 sky130_fd_sc_hd__xnor2_2 _19909_ (.A(_01729_),
    .B(_01730_),
    .Y(_01731_));
 sky130_fd_sc_hd__xnor2_2 _19910_ (.A(_01718_),
    .B(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__a21oi_1 _19911_ (.A1(_01717_),
    .A2(_01732_),
    .B1(_07576_),
    .Y(_01733_));
 sky130_fd_sc_hd__o21ai_2 _19912_ (.A1(_01717_),
    .A2(_01732_),
    .B1(_01733_),
    .Y(_01734_));
 sky130_fd_sc_hd__o211a_1 _19913_ (.A1(net907),
    .A2(_10616_),
    .B1(_01734_),
    .C1(_11714_),
    .X(_00745_));
 sky130_fd_sc_hd__buf_4 _19914_ (.A(_05787_),
    .X(_01735_));
 sky130_fd_sc_hd__and2b_1 _19915_ (.A_N(_01729_),
    .B(_01730_),
    .X(_01736_));
 sky130_fd_sc_hd__a21o_1 _19916_ (.A1(_01721_),
    .A2(_01724_),
    .B1(_01723_),
    .X(_01737_));
 sky130_fd_sc_hd__a21o_2 _19917_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[19] ),
    .A2(_01395_),
    .B1(_01396_),
    .X(_01738_));
 sky130_fd_sc_hd__xnor2_1 _19918_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[20] ),
    .B(_01480_),
    .Y(_01739_));
 sky130_fd_sc_hd__nor2_1 _19919_ (.A(_01561_),
    .B(_01739_),
    .Y(_01740_));
 sky130_fd_sc_hd__and2_1 _19920_ (.A(_01561_),
    .B(_01739_),
    .X(_01741_));
 sky130_fd_sc_hd__nor2_2 _19921_ (.A(_01740_),
    .B(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__xor2_4 _19922_ (.A(_01738_),
    .B(_01742_),
    .X(_01743_));
 sky130_fd_sc_hd__nor2_1 _19923_ (.A(_01611_),
    .B(_01726_),
    .Y(_01744_));
 sky130_fd_sc_hd__xor2_2 _19924_ (.A(_01743_),
    .B(_01744_),
    .X(_01745_));
 sky130_fd_sc_hd__xnor2_1 _19925_ (.A(_01737_),
    .B(_01745_),
    .Y(_01746_));
 sky130_fd_sc_hd__a22o_1 _19926_ (.A1(_01720_),
    .A2(_01728_),
    .B1(_01744_),
    .B2(_01701_),
    .X(_01747_));
 sky130_fd_sc_hd__xnor2_1 _19927_ (.A(_01746_),
    .B(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__xor2_1 _19928_ (.A(_01736_),
    .B(_01748_),
    .X(_01749_));
 sky130_fd_sc_hd__and2_1 _19929_ (.A(_01709_),
    .B(_01732_),
    .X(_01750_));
 sky130_fd_sc_hd__and3_1 _19930_ (.A(_01673_),
    .B(_01694_),
    .C(_01750_),
    .X(_01751_));
 sky130_fd_sc_hd__nand2_1 _19931_ (.A(_01718_),
    .B(_01716_),
    .Y(_01752_));
 sky130_fd_sc_hd__a22o_1 _19932_ (.A1(_01710_),
    .A2(_01750_),
    .B1(_01752_),
    .B2(_01731_),
    .X(_01753_));
 sky130_fd_sc_hd__a21o_1 _19933_ (.A1(_01652_),
    .A2(_01751_),
    .B1(_01753_),
    .X(_01754_));
 sky130_fd_sc_hd__nand2_1 _19934_ (.A(_01749_),
    .B(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hd__or2_1 _19935_ (.A(_01749_),
    .B(_01754_),
    .X(_01756_));
 sky130_fd_sc_hd__a21o_1 _19936_ (.A1(_01755_),
    .A2(_01756_),
    .B1(_06682_),
    .X(_01757_));
 sky130_fd_sc_hd__o211a_1 _19937_ (.A1(net925),
    .A2(_01735_),
    .B1(_01757_),
    .C1(_11714_),
    .X(_00746_));
 sky130_fd_sc_hd__nand2_1 _19938_ (.A(_01736_),
    .B(_01748_),
    .Y(_01758_));
 sky130_fd_sc_hd__or2b_1 _19939_ (.A(_01746_),
    .B_N(_01747_),
    .X(_01759_));
 sky130_fd_sc_hd__a21o_1 _19940_ (.A1(_01738_),
    .A2(_01742_),
    .B1(_01740_),
    .X(_01760_));
 sky130_fd_sc_hd__buf_2 _19941_ (.A(_01395_),
    .X(_01761_));
 sky130_fd_sc_hd__clkbuf_4 _19942_ (.A(_01396_),
    .X(_01762_));
 sky130_fd_sc_hd__a21o_1 _19943_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[20] ),
    .A2(_01761_),
    .B1(_01762_),
    .X(_01763_));
 sky130_fd_sc_hd__buf_4 _19944_ (.A(_01480_),
    .X(_01764_));
 sky130_fd_sc_hd__xnor2_1 _19945_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[21] ),
    .B(_01764_),
    .Y(_01765_));
 sky130_fd_sc_hd__nor2_1 _19946_ (.A(_01561_),
    .B(_01765_),
    .Y(_01766_));
 sky130_fd_sc_hd__and2_1 _19947_ (.A(_01561_),
    .B(_01765_),
    .X(_01767_));
 sky130_fd_sc_hd__nor2_1 _19948_ (.A(_01766_),
    .B(_01767_),
    .Y(_01768_));
 sky130_fd_sc_hd__xor2_2 _19949_ (.A(_01763_),
    .B(_01768_),
    .X(_01769_));
 sky130_fd_sc_hd__nor2_2 _19950_ (.A(_01611_),
    .B(_01743_),
    .Y(_01770_));
 sky130_fd_sc_hd__xor2_2 _19951_ (.A(_01769_),
    .B(_01770_),
    .X(_01771_));
 sky130_fd_sc_hd__xnor2_2 _19952_ (.A(_01760_),
    .B(_01771_),
    .Y(_01772_));
 sky130_fd_sc_hd__a22oi_4 _19953_ (.A1(_01737_),
    .A2(_01745_),
    .B1(_01770_),
    .B2(_01726_),
    .Y(_01773_));
 sky130_fd_sc_hd__xor2_1 _19954_ (.A(_01772_),
    .B(_01773_),
    .X(_01774_));
 sky130_fd_sc_hd__xnor2_1 _19955_ (.A(_01759_),
    .B(_01774_),
    .Y(_01775_));
 sky130_fd_sc_hd__a21oi_1 _19956_ (.A1(_01758_),
    .A2(_01755_),
    .B1(_01775_),
    .Y(_01776_));
 sky130_fd_sc_hd__a31o_1 _19957_ (.A1(_01758_),
    .A2(_01755_),
    .A3(_01775_),
    .B1(_10957_),
    .X(_01777_));
 sky130_fd_sc_hd__o221a_1 _19958_ (.A1(net1095),
    .A2(_01202_),
    .B1(_01776_),
    .B2(_01777_),
    .C1(_11228_),
    .X(_00747_));
 sky130_fd_sc_hd__a21o_1 _19959_ (.A1(_01763_),
    .A2(_01768_),
    .B1(_01766_),
    .X(_01778_));
 sky130_fd_sc_hd__a21o_1 _19960_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[21] ),
    .A2(_01761_),
    .B1(_01762_),
    .X(_01779_));
 sky130_fd_sc_hd__xnor2_2 _19961_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[22] ),
    .B(_01764_),
    .Y(_01780_));
 sky130_fd_sc_hd__xor2_2 _19962_ (.A(_01561_),
    .B(_01780_),
    .X(_01781_));
 sky130_fd_sc_hd__xor2_2 _19963_ (.A(_01779_),
    .B(_01781_),
    .X(_01782_));
 sky130_fd_sc_hd__clkbuf_4 _19964_ (.A(_01611_),
    .X(_01783_));
 sky130_fd_sc_hd__nor2_1 _19965_ (.A(_01783_),
    .B(_01769_),
    .Y(_01784_));
 sky130_fd_sc_hd__xor2_2 _19966_ (.A(_01782_),
    .B(_01784_),
    .X(_01785_));
 sky130_fd_sc_hd__xnor2_1 _19967_ (.A(_01778_),
    .B(_01785_),
    .Y(_01786_));
 sky130_fd_sc_hd__a22oi_2 _19968_ (.A1(_01760_),
    .A2(_01771_),
    .B1(_01784_),
    .B2(_01743_),
    .Y(_01787_));
 sky130_fd_sc_hd__nor2_1 _19969_ (.A(_01786_),
    .B(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__and2_1 _19970_ (.A(_01786_),
    .B(_01787_),
    .X(_01789_));
 sky130_fd_sc_hd__nor4_1 _19971_ (.A(_01772_),
    .B(_01773_),
    .C(_01788_),
    .D(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__o22a_1 _19972_ (.A1(_01772_),
    .A2(_01773_),
    .B1(_01788_),
    .B2(_01789_),
    .X(_01791_));
 sky130_fd_sc_hd__nor2_1 _19973_ (.A(_01790_),
    .B(_01791_),
    .Y(_01792_));
 sky130_fd_sc_hd__and2_1 _19974_ (.A(_01749_),
    .B(_01775_),
    .X(_01793_));
 sky130_fd_sc_hd__a21boi_1 _19975_ (.A1(_01759_),
    .A2(_01758_),
    .B1_N(_01774_),
    .Y(_01794_));
 sky130_fd_sc_hd__a21o_1 _19976_ (.A1(_01754_),
    .A2(_01793_),
    .B1(_01794_),
    .X(_01795_));
 sky130_fd_sc_hd__xor2_2 _19977_ (.A(_01792_),
    .B(_01795_),
    .X(_01796_));
 sky130_fd_sc_hd__or2_1 _19978_ (.A(net825),
    .B(_01386_),
    .X(_01797_));
 sky130_fd_sc_hd__o211a_1 _19979_ (.A1(_11177_),
    .A2(_01796_),
    .B1(_01797_),
    .C1(_11714_),
    .X(_00748_));
 sky130_fd_sc_hd__a21oi_1 _19980_ (.A1(_01792_),
    .A2(_01795_),
    .B1(net168),
    .Y(_01798_));
 sky130_fd_sc_hd__nor2_1 _19981_ (.A(_01563_),
    .B(_01780_),
    .Y(_01799_));
 sky130_fd_sc_hd__a21o_1 _19982_ (.A1(_01779_),
    .A2(_01781_),
    .B1(_01799_),
    .X(_01800_));
 sky130_fd_sc_hd__a21o_1 _19983_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[22] ),
    .A2(_01761_),
    .B1(_01762_),
    .X(_01801_));
 sky130_fd_sc_hd__xnor2_1 _19984_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[23] ),
    .B(_01764_),
    .Y(_01802_));
 sky130_fd_sc_hd__nor2_1 _19985_ (.A(_01561_),
    .B(_01802_),
    .Y(_01803_));
 sky130_fd_sc_hd__nand2_1 _19986_ (.A(_01561_),
    .B(_01802_),
    .Y(_01804_));
 sky130_fd_sc_hd__and2b_1 _19987_ (.A_N(_01803_),
    .B(_01804_),
    .X(_01805_));
 sky130_fd_sc_hd__xor2_2 _19988_ (.A(_01801_),
    .B(_01805_),
    .X(_01806_));
 sky130_fd_sc_hd__nor2_1 _19989_ (.A(_01783_),
    .B(_01782_),
    .Y(_01807_));
 sky130_fd_sc_hd__xor2_1 _19990_ (.A(_01806_),
    .B(_01807_),
    .X(_01808_));
 sky130_fd_sc_hd__nand2_1 _19991_ (.A(_01800_),
    .B(_01808_),
    .Y(_01809_));
 sky130_fd_sc_hd__or2_1 _19992_ (.A(_01800_),
    .B(_01808_),
    .X(_01810_));
 sky130_fd_sc_hd__nand2_1 _19993_ (.A(_01809_),
    .B(_01810_),
    .Y(_01811_));
 sky130_fd_sc_hd__a22oi_2 _19994_ (.A1(_01778_),
    .A2(_01785_),
    .B1(_01807_),
    .B2(_01769_),
    .Y(_01812_));
 sky130_fd_sc_hd__nor2_2 _19995_ (.A(_01811_),
    .B(_01812_),
    .Y(_01813_));
 sky130_fd_sc_hd__and2_1 _19996_ (.A(_01811_),
    .B(_01812_),
    .X(_01814_));
 sky130_fd_sc_hd__nor2_1 _19997_ (.A(_01813_),
    .B(_01814_),
    .Y(_01815_));
 sky130_fd_sc_hd__xor2_1 _19998_ (.A(_01788_),
    .B(_01815_),
    .X(_01816_));
 sky130_fd_sc_hd__nor2_1 _19999_ (.A(_01798_),
    .B(_01816_),
    .Y(_01817_));
 sky130_fd_sc_hd__a21o_1 _20000_ (.A1(_01798_),
    .A2(_01816_),
    .B1(_09292_),
    .X(_01818_));
 sky130_fd_sc_hd__o221a_1 _20001_ (.A1(net1094),
    .A2(_01202_),
    .B1(_01817_),
    .B2(_01818_),
    .C1(_11228_),
    .X(_00749_));
 sky130_fd_sc_hd__buf_4 _20002_ (.A(_07057_),
    .X(_01819_));
 sky130_fd_sc_hd__and2_1 _20003_ (.A(_01792_),
    .B(_01816_),
    .X(_01820_));
 sky130_fd_sc_hd__or2_1 _20004_ (.A(_01788_),
    .B(net168),
    .X(_01821_));
 sky130_fd_sc_hd__a21o_1 _20005_ (.A1(_01753_),
    .A2(_01793_),
    .B1(_01794_),
    .X(_01822_));
 sky130_fd_sc_hd__a22o_1 _20006_ (.A1(_01815_),
    .A2(_01821_),
    .B1(_01822_),
    .B2(_01820_),
    .X(_01823_));
 sky130_fd_sc_hd__a41o_4 _20007_ (.A1(_01652_),
    .A2(_01751_),
    .A3(_01793_),
    .A4(_01820_),
    .B1(_01823_),
    .X(_01824_));
 sky130_fd_sc_hd__nor2_1 _20008_ (.A(_01783_),
    .B(_01806_),
    .Y(_01825_));
 sky130_fd_sc_hd__nand2_1 _20009_ (.A(_01782_),
    .B(_01825_),
    .Y(_01826_));
 sky130_fd_sc_hd__a21o_1 _20010_ (.A1(_01801_),
    .A2(_01804_),
    .B1(_01803_),
    .X(_01827_));
 sky130_fd_sc_hd__a21o_1 _20011_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[23] ),
    .A2(_01761_),
    .B1(_01762_),
    .X(_01828_));
 sky130_fd_sc_hd__xnor2_2 _20012_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[24] ),
    .B(_01764_),
    .Y(_01829_));
 sky130_fd_sc_hd__xor2_2 _20013_ (.A(_01561_),
    .B(_01829_),
    .X(_01830_));
 sky130_fd_sc_hd__xor2_2 _20014_ (.A(_01828_),
    .B(_01830_),
    .X(_01831_));
 sky130_fd_sc_hd__xor2_1 _20015_ (.A(_01831_),
    .B(_01825_),
    .X(_01832_));
 sky130_fd_sc_hd__xnor2_1 _20016_ (.A(_01827_),
    .B(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__a21o_1 _20017_ (.A1(_01809_),
    .A2(_01826_),
    .B1(_01833_),
    .X(_01834_));
 sky130_fd_sc_hd__nand3_1 _20018_ (.A(_01809_),
    .B(_01833_),
    .C(_01826_),
    .Y(_01835_));
 sky130_fd_sc_hd__and2_1 _20019_ (.A(_01834_),
    .B(_01835_),
    .X(_01836_));
 sky130_fd_sc_hd__xor2_2 _20020_ (.A(_01813_),
    .B(_01836_),
    .X(_01837_));
 sky130_fd_sc_hd__xor2_2 _20021_ (.A(_01824_),
    .B(_01837_),
    .X(_01838_));
 sky130_fd_sc_hd__or2_1 _20022_ (.A(net786),
    .B(_01386_),
    .X(_01839_));
 sky130_fd_sc_hd__clkbuf_4 _20023_ (.A(_10447_),
    .X(_01840_));
 sky130_fd_sc_hd__o211a_1 _20024_ (.A1(_01819_),
    .A2(_01838_),
    .B1(_01839_),
    .C1(_01840_),
    .X(_00750_));
 sky130_fd_sc_hd__nand2_1 _20025_ (.A(_01813_),
    .B(_01836_),
    .Y(_01841_));
 sky130_fd_sc_hd__nand2_1 _20026_ (.A(_01824_),
    .B(_01837_),
    .Y(_01842_));
 sky130_fd_sc_hd__nor2_1 _20027_ (.A(_01563_),
    .B(_01829_),
    .Y(_01843_));
 sky130_fd_sc_hd__a21o_1 _20028_ (.A1(_01828_),
    .A2(_01830_),
    .B1(_01843_),
    .X(_01844_));
 sky130_fd_sc_hd__a21o_1 _20029_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[24] ),
    .A2(_01761_),
    .B1(_01762_),
    .X(_01845_));
 sky130_fd_sc_hd__xnor2_1 _20030_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[25] ),
    .B(_01764_),
    .Y(_01846_));
 sky130_fd_sc_hd__nor2_1 _20031_ (.A(_01561_),
    .B(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__nand2_1 _20032_ (.A(_01562_),
    .B(_01846_),
    .Y(_01848_));
 sky130_fd_sc_hd__and2b_1 _20033_ (.A_N(_01847_),
    .B(_01848_),
    .X(_01849_));
 sky130_fd_sc_hd__xor2_2 _20034_ (.A(_01845_),
    .B(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__nor2_1 _20035_ (.A(_01783_),
    .B(_01831_),
    .Y(_01851_));
 sky130_fd_sc_hd__xor2_1 _20036_ (.A(_01850_),
    .B(_01851_),
    .X(_01852_));
 sky130_fd_sc_hd__nand2_1 _20037_ (.A(_01844_),
    .B(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__or2_1 _20038_ (.A(_01844_),
    .B(_01852_),
    .X(_01854_));
 sky130_fd_sc_hd__nand2_1 _20039_ (.A(_01853_),
    .B(_01854_),
    .Y(_01855_));
 sky130_fd_sc_hd__a22oi_1 _20040_ (.A1(_01827_),
    .A2(_01832_),
    .B1(_01851_),
    .B2(_01806_),
    .Y(_01856_));
 sky130_fd_sc_hd__nor2_1 _20041_ (.A(_01855_),
    .B(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__and2_1 _20042_ (.A(_01855_),
    .B(_01856_),
    .X(_01858_));
 sky130_fd_sc_hd__nor2_1 _20043_ (.A(_01857_),
    .B(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__xnor2_1 _20044_ (.A(_01834_),
    .B(_01859_),
    .Y(_01860_));
 sky130_fd_sc_hd__a21oi_1 _20045_ (.A1(_01841_),
    .A2(_01842_),
    .B1(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hd__a31o_1 _20046_ (.A1(_01841_),
    .A2(_01842_),
    .A3(_01860_),
    .B1(_10957_),
    .X(_01862_));
 sky130_fd_sc_hd__clkbuf_8 _20047_ (.A(_07707_),
    .X(_01863_));
 sky130_fd_sc_hd__o221a_1 _20048_ (.A1(net1099),
    .A2(_01202_),
    .B1(_01861_),
    .B2(_01862_),
    .C1(_01863_),
    .X(_00751_));
 sky130_fd_sc_hd__a21boi_2 _20049_ (.A1(_01834_),
    .A2(_01841_),
    .B1_N(_01859_),
    .Y(_01864_));
 sky130_fd_sc_hd__nand2_1 _20050_ (.A(_01837_),
    .B(_01860_),
    .Y(_01865_));
 sky130_fd_sc_hd__inv_2 _20051_ (.A(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__and2_1 _20052_ (.A(_01824_),
    .B(_01866_),
    .X(_01867_));
 sky130_fd_sc_hd__nor2_1 _20053_ (.A(_01783_),
    .B(_01850_),
    .Y(_01868_));
 sky130_fd_sc_hd__nand2_1 _20054_ (.A(_01831_),
    .B(_01868_),
    .Y(_01869_));
 sky130_fd_sc_hd__a21o_1 _20055_ (.A1(_01845_),
    .A2(_01848_),
    .B1(_01847_),
    .X(_01870_));
 sky130_fd_sc_hd__a21o_1 _20056_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[25] ),
    .A2(_01761_),
    .B1(_01762_),
    .X(_01871_));
 sky130_fd_sc_hd__xnor2_1 _20057_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[26] ),
    .B(_01764_),
    .Y(_01872_));
 sky130_fd_sc_hd__nor2_1 _20058_ (.A(_01562_),
    .B(_01872_),
    .Y(_01873_));
 sky130_fd_sc_hd__nand2_1 _20059_ (.A(_01562_),
    .B(_01872_),
    .Y(_01874_));
 sky130_fd_sc_hd__and2b_1 _20060_ (.A_N(_01873_),
    .B(_01874_),
    .X(_01875_));
 sky130_fd_sc_hd__xor2_2 _20061_ (.A(_01871_),
    .B(_01875_),
    .X(_01876_));
 sky130_fd_sc_hd__xor2_2 _20062_ (.A(_01876_),
    .B(_01868_),
    .X(_01877_));
 sky130_fd_sc_hd__xnor2_1 _20063_ (.A(_01870_),
    .B(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__a21o_1 _20064_ (.A1(_01853_),
    .A2(_01869_),
    .B1(_01878_),
    .X(_01879_));
 sky130_fd_sc_hd__nand3_1 _20065_ (.A(_01853_),
    .B(_01878_),
    .C(_01869_),
    .Y(_01880_));
 sky130_fd_sc_hd__and2_1 _20066_ (.A(_01879_),
    .B(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__nand2_1 _20067_ (.A(_01857_),
    .B(_01881_),
    .Y(_01882_));
 sky130_fd_sc_hd__or2_1 _20068_ (.A(_01857_),
    .B(_01881_),
    .X(_01883_));
 sky130_fd_sc_hd__and2_1 _20069_ (.A(_01882_),
    .B(_01883_),
    .X(_01884_));
 sky130_fd_sc_hd__o21ai_2 _20070_ (.A1(_01864_),
    .A2(_01867_),
    .B1(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__or3_1 _20071_ (.A(_01884_),
    .B(_01864_),
    .C(_01867_),
    .X(_01886_));
 sky130_fd_sc_hd__and2_1 _20072_ (.A(\top_inst.deskew_buff_inst.col_input[26] ),
    .B(_05730_),
    .X(_01887_));
 sky130_fd_sc_hd__a31o_1 _20073_ (.A1(_05887_),
    .A2(_01885_),
    .A3(_01886_),
    .B1(_01887_),
    .X(_01888_));
 sky130_fd_sc_hd__and2_1 _20074_ (.A(_11722_),
    .B(_01888_),
    .X(_01889_));
 sky130_fd_sc_hd__clkbuf_1 _20075_ (.A(_01889_),
    .X(_00752_));
 sky130_fd_sc_hd__a21o_1 _20076_ (.A1(_01871_),
    .A2(_01874_),
    .B1(_01873_),
    .X(_01890_));
 sky130_fd_sc_hd__a21o_2 _20077_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[26] ),
    .A2(_01761_),
    .B1(_01762_),
    .X(_01891_));
 sky130_fd_sc_hd__xnor2_1 _20078_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[27] ),
    .B(_01764_),
    .Y(_01892_));
 sky130_fd_sc_hd__nor2_1 _20079_ (.A(_01562_),
    .B(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hd__nand2_1 _20080_ (.A(_01562_),
    .B(_01892_),
    .Y(_01894_));
 sky130_fd_sc_hd__and2b_1 _20081_ (.A_N(_01893_),
    .B(_01894_),
    .X(_01895_));
 sky130_fd_sc_hd__xor2_4 _20082_ (.A(_01891_),
    .B(_01895_),
    .X(_01896_));
 sky130_fd_sc_hd__nor2_1 _20083_ (.A(_01783_),
    .B(_01876_),
    .Y(_01897_));
 sky130_fd_sc_hd__xor2_1 _20084_ (.A(_01896_),
    .B(_01897_),
    .X(_01898_));
 sky130_fd_sc_hd__nand2_1 _20085_ (.A(_01890_),
    .B(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__or2_1 _20086_ (.A(_01890_),
    .B(_01898_),
    .X(_01900_));
 sky130_fd_sc_hd__nand2_1 _20087_ (.A(_01899_),
    .B(_01900_),
    .Y(_01901_));
 sky130_fd_sc_hd__a22oi_2 _20088_ (.A1(_01870_),
    .A2(_01877_),
    .B1(_01897_),
    .B2(_01850_),
    .Y(_01902_));
 sky130_fd_sc_hd__nor2_1 _20089_ (.A(_01901_),
    .B(_01902_),
    .Y(_01903_));
 sky130_fd_sc_hd__and2_1 _20090_ (.A(_01901_),
    .B(_01902_),
    .X(_01904_));
 sky130_fd_sc_hd__nor2_1 _20091_ (.A(_01903_),
    .B(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__xnor2_2 _20092_ (.A(_01879_),
    .B(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hd__a21oi_1 _20093_ (.A1(_01882_),
    .A2(_01885_),
    .B1(_01906_),
    .Y(_01907_));
 sky130_fd_sc_hd__a31o_1 _20094_ (.A1(_01882_),
    .A2(_01885_),
    .A3(_01906_),
    .B1(_10957_),
    .X(_01908_));
 sky130_fd_sc_hd__o221a_1 _20095_ (.A1(net1098),
    .A2(_01202_),
    .B1(_01907_),
    .B2(_01908_),
    .C1(_01863_),
    .X(_00753_));
 sky130_fd_sc_hd__and3_1 _20096_ (.A(_01884_),
    .B(_01866_),
    .C(_01906_),
    .X(_01909_));
 sky130_fd_sc_hd__nand2_1 _20097_ (.A(_01879_),
    .B(_01882_),
    .Y(_01910_));
 sky130_fd_sc_hd__a32o_1 _20098_ (.A1(_01884_),
    .A2(_01864_),
    .A3(_01906_),
    .B1(_01910_),
    .B2(_01905_),
    .X(_01911_));
 sky130_fd_sc_hd__a21o_1 _20099_ (.A1(_01824_),
    .A2(_01909_),
    .B1(_01911_),
    .X(_01912_));
 sky130_fd_sc_hd__nor2_1 _20100_ (.A(_01783_),
    .B(_01896_),
    .Y(_01913_));
 sky130_fd_sc_hd__nand2_1 _20101_ (.A(_01876_),
    .B(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__a21o_1 _20102_ (.A1(_01891_),
    .A2(_01894_),
    .B1(_01893_),
    .X(_01915_));
 sky130_fd_sc_hd__a21o_1 _20103_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[27] ),
    .A2(_01761_),
    .B1(_01762_),
    .X(_01916_));
 sky130_fd_sc_hd__xnor2_1 _20104_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[28] ),
    .B(_01764_),
    .Y(_01917_));
 sky130_fd_sc_hd__or2_1 _20105_ (.A(_01563_),
    .B(_01917_),
    .X(_01918_));
 sky130_fd_sc_hd__nand2_1 _20106_ (.A(_01563_),
    .B(_01917_),
    .Y(_01919_));
 sky130_fd_sc_hd__and2_1 _20107_ (.A(_01918_),
    .B(_01919_),
    .X(_01920_));
 sky130_fd_sc_hd__xor2_2 _20108_ (.A(_01916_),
    .B(_01920_),
    .X(_01921_));
 sky130_fd_sc_hd__xor2_2 _20109_ (.A(_01921_),
    .B(_01913_),
    .X(_01922_));
 sky130_fd_sc_hd__xnor2_1 _20110_ (.A(_01915_),
    .B(_01922_),
    .Y(_01923_));
 sky130_fd_sc_hd__a21o_1 _20111_ (.A1(_01899_),
    .A2(_01914_),
    .B1(_01923_),
    .X(_01924_));
 sky130_fd_sc_hd__nand3_1 _20112_ (.A(_01899_),
    .B(_01923_),
    .C(_01914_),
    .Y(_01925_));
 sky130_fd_sc_hd__and2_1 _20113_ (.A(_01924_),
    .B(_01925_),
    .X(_01926_));
 sky130_fd_sc_hd__nand2_1 _20114_ (.A(_01903_),
    .B(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__or2_1 _20115_ (.A(_01903_),
    .B(_01926_),
    .X(_01928_));
 sky130_fd_sc_hd__and2_1 _20116_ (.A(_01927_),
    .B(_01928_),
    .X(_01929_));
 sky130_fd_sc_hd__xor2_2 _20117_ (.A(_01912_),
    .B(_01929_),
    .X(_01930_));
 sky130_fd_sc_hd__or2_1 _20118_ (.A(net756),
    .B(_01386_),
    .X(_01931_));
 sky130_fd_sc_hd__o211a_1 _20119_ (.A1(_01819_),
    .A2(_01930_),
    .B1(_01931_),
    .C1(_01840_),
    .X(_00754_));
 sky130_fd_sc_hd__a21boi_1 _20120_ (.A1(_01912_),
    .A2(_01929_),
    .B1_N(_01927_),
    .Y(_01932_));
 sky130_fd_sc_hd__nand2_1 _20121_ (.A(_01916_),
    .B(_01920_),
    .Y(_01933_));
 sky130_fd_sc_hd__a21o_1 _20122_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[28] ),
    .A2(_01761_),
    .B1(_01762_),
    .X(_01934_));
 sky130_fd_sc_hd__xnor2_1 _20123_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[29] ),
    .B(_01764_),
    .Y(_01935_));
 sky130_fd_sc_hd__nor2_1 _20124_ (.A(_01563_),
    .B(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__nand2_1 _20125_ (.A(_01563_),
    .B(_01935_),
    .Y(_01937_));
 sky130_fd_sc_hd__and2b_1 _20126_ (.A_N(_01936_),
    .B(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__xor2_2 _20127_ (.A(_01934_),
    .B(_01938_),
    .X(_01939_));
 sky130_fd_sc_hd__nor2_2 _20128_ (.A(_01783_),
    .B(_01921_),
    .Y(_01940_));
 sky130_fd_sc_hd__xnor2_1 _20129_ (.A(_01939_),
    .B(_01940_),
    .Y(_01941_));
 sky130_fd_sc_hd__a21oi_1 _20130_ (.A1(_01918_),
    .A2(_01933_),
    .B1(_01941_),
    .Y(_01942_));
 sky130_fd_sc_hd__and3_1 _20131_ (.A(_01918_),
    .B(_01933_),
    .C(_01941_),
    .X(_01943_));
 sky130_fd_sc_hd__or2_1 _20132_ (.A(_01942_),
    .B(_01943_),
    .X(_01944_));
 sky130_fd_sc_hd__a22oi_4 _20133_ (.A1(_01915_),
    .A2(_01922_),
    .B1(_01940_),
    .B2(_01896_),
    .Y(_01945_));
 sky130_fd_sc_hd__xor2_1 _20134_ (.A(_01944_),
    .B(_01945_),
    .X(_01946_));
 sky130_fd_sc_hd__xnor2_1 _20135_ (.A(_01924_),
    .B(_01946_),
    .Y(_01947_));
 sky130_fd_sc_hd__o21ai_1 _20136_ (.A1(_01932_),
    .A2(_01947_),
    .B1(_05316_),
    .Y(_01948_));
 sky130_fd_sc_hd__a21o_1 _20137_ (.A1(_01932_),
    .A2(_01947_),
    .B1(_01948_),
    .X(_01949_));
 sky130_fd_sc_hd__o211a_1 _20138_ (.A1(net790),
    .A2(_01735_),
    .B1(_01949_),
    .C1(_01840_),
    .X(_00755_));
 sky130_fd_sc_hd__a21o_1 _20139_ (.A1(_01934_),
    .A2(_01937_),
    .B1(_01936_),
    .X(_01950_));
 sky130_fd_sc_hd__a21o_1 _20140_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[29] ),
    .A2(_01761_),
    .B1(_01762_),
    .X(_01951_));
 sky130_fd_sc_hd__xnor2_1 _20141_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[30] ),
    .B(_01764_),
    .Y(_01952_));
 sky130_fd_sc_hd__nor2_1 _20142_ (.A(_01563_),
    .B(_01952_),
    .Y(_01953_));
 sky130_fd_sc_hd__and2_1 _20143_ (.A(_01563_),
    .B(_01952_),
    .X(_01954_));
 sky130_fd_sc_hd__nor2_1 _20144_ (.A(_01953_),
    .B(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__xor2_1 _20145_ (.A(_01951_),
    .B(_01955_),
    .X(_01956_));
 sky130_fd_sc_hd__nor2_1 _20146_ (.A(_01783_),
    .B(_01939_),
    .Y(_01957_));
 sky130_fd_sc_hd__xor2_1 _20147_ (.A(_01956_),
    .B(_01957_),
    .X(_01958_));
 sky130_fd_sc_hd__xnor2_1 _20148_ (.A(_01950_),
    .B(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__a21oi_1 _20149_ (.A1(_01921_),
    .A2(_01957_),
    .B1(_01942_),
    .Y(_01960_));
 sky130_fd_sc_hd__or2_1 _20150_ (.A(_01959_),
    .B(_01960_),
    .X(_01961_));
 sky130_fd_sc_hd__nand2_1 _20151_ (.A(_01959_),
    .B(_01960_),
    .Y(_01962_));
 sky130_fd_sc_hd__and2_1 _20152_ (.A(_01961_),
    .B(_01962_),
    .X(_01963_));
 sky130_fd_sc_hd__or3b_1 _20153_ (.A(_01944_),
    .B(_01945_),
    .C_N(_01963_),
    .X(_01964_));
 sky130_fd_sc_hd__o21bai_1 _20154_ (.A1(_01944_),
    .A2(_01945_),
    .B1_N(_01963_),
    .Y(_01965_));
 sky130_fd_sc_hd__and2_1 _20155_ (.A(_01964_),
    .B(_01965_),
    .X(_01966_));
 sky130_fd_sc_hd__nand2_1 _20156_ (.A(_01924_),
    .B(_01927_),
    .Y(_01967_));
 sky130_fd_sc_hd__a32o_2 _20157_ (.A1(_01912_),
    .A2(_01929_),
    .A3(_01947_),
    .B1(_01967_),
    .B2(_01946_),
    .X(_01968_));
 sky130_fd_sc_hd__nand2_2 _20158_ (.A(_01968_),
    .B(_01966_),
    .Y(_01969_));
 sky130_fd_sc_hd__o21a_1 _20159_ (.A1(_01966_),
    .A2(_01968_),
    .B1(_10831_),
    .X(_01970_));
 sky130_fd_sc_hd__a22o_1 _20160_ (.A1(\top_inst.deskew_buff_inst.col_input[30] ),
    .A2(_11723_),
    .B1(_01969_),
    .B2(_01970_),
    .X(_01971_));
 sky130_fd_sc_hd__and2_4 _20161_ (.A(_11722_),
    .B(_01971_),
    .X(_01972_));
 sky130_fd_sc_hd__clkbuf_1 _20162_ (.A(_01972_),
    .X(_00756_));
 sky130_fd_sc_hd__a21oi_1 _20163_ (.A1(_01951_),
    .A2(_01955_),
    .B1(_01953_),
    .Y(_01973_));
 sky130_fd_sc_hd__xnor2_1 _20164_ (.A(_01961_),
    .B(_01973_),
    .Y(_01974_));
 sky130_fd_sc_hd__o21a_1 _20165_ (.A1(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[30] ),
    .A2(_01352_),
    .B1(_01524_),
    .X(_01975_));
 sky130_fd_sc_hd__nor2_1 _20166_ (.A(_01783_),
    .B(_01956_),
    .Y(_01976_));
 sky130_fd_sc_hd__a22o_1 _20167_ (.A1(_01950_),
    .A2(_01958_),
    .B1(_01976_),
    .B2(_01939_),
    .X(_01977_));
 sky130_fd_sc_hd__xnor2_1 _20168_ (.A(_01563_),
    .B(_01977_),
    .Y(_01978_));
 sky130_fd_sc_hd__xnor2_1 _20169_ (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[31] ),
    .B(_01976_),
    .Y(_01979_));
 sky130_fd_sc_hd__xnor2_1 _20170_ (.A(_01978_),
    .B(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__xnor2_1 _20171_ (.A(_01975_),
    .B(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__xnor2_2 _20172_ (.A(_01974_),
    .B(_01981_),
    .Y(_01982_));
 sky130_fd_sc_hd__a21oi_1 _20173_ (.A1(_01964_),
    .A2(_01969_),
    .B1(_01982_),
    .Y(_01983_));
 sky130_fd_sc_hd__buf_8 _20174_ (.A(_05633_),
    .X(_01984_));
 sky130_fd_sc_hd__a31o_1 _20175_ (.A1(_01964_),
    .A2(_01969_),
    .A3(_01982_),
    .B1(_01984_),
    .X(_01985_));
 sky130_fd_sc_hd__o221a_1 _20176_ (.A1(net490),
    .A2(_01202_),
    .B1(_01983_),
    .B2(_01985_),
    .C1(_01863_),
    .X(_00757_));
 sky130_fd_sc_hd__buf_2 _20177_ (.A(\top_inst.grid_inst.data_path_wires[16][0] ),
    .X(_01986_));
 sky130_fd_sc_hd__clkbuf_4 _20178_ (.A(_01986_),
    .X(_01987_));
 sky130_fd_sc_hd__or2_1 _20179_ (.A(_10030_),
    .B(_11677_),
    .X(_01988_));
 sky130_fd_sc_hd__o211a_1 _20180_ (.A1(_01987_),
    .A2(_10033_),
    .B1(_01988_),
    .C1(_01840_),
    .X(_00758_));
 sky130_fd_sc_hd__clkbuf_4 _20181_ (.A(\top_inst.grid_inst.data_path_wires[16][1] ),
    .X(_01989_));
 sky130_fd_sc_hd__buf_4 _20182_ (.A(_01989_),
    .X(_01990_));
 sky130_fd_sc_hd__or2_1 _20183_ (.A(_10030_),
    .B(_11682_),
    .X(_01991_));
 sky130_fd_sc_hd__o211a_1 _20184_ (.A1(_01990_),
    .A2(_10033_),
    .B1(_01991_),
    .C1(_01840_),
    .X(_00759_));
 sky130_fd_sc_hd__buf_2 _20185_ (.A(\top_inst.grid_inst.data_path_wires[16][2] ),
    .X(_01992_));
 sky130_fd_sc_hd__buf_4 _20186_ (.A(_01992_),
    .X(_01993_));
 sky130_fd_sc_hd__or2_2 _20187_ (.A(_10030_),
    .B(_11687_),
    .X(_01994_));
 sky130_fd_sc_hd__o211a_1 _20188_ (.A1(_01993_),
    .A2(_10033_),
    .B1(_01994_),
    .C1(_01840_),
    .X(_00760_));
 sky130_fd_sc_hd__buf_4 _20189_ (.A(\top_inst.grid_inst.data_path_wires[16][3] ),
    .X(_01995_));
 sky130_fd_sc_hd__or2_2 _20190_ (.A(_10030_),
    .B(_11692_),
    .X(_01996_));
 sky130_fd_sc_hd__o211a_1 _20191_ (.A1(_01995_),
    .A2(_10033_),
    .B1(_01996_),
    .C1(_01840_),
    .X(_00761_));
 sky130_fd_sc_hd__buf_4 _20192_ (.A(\top_inst.grid_inst.data_path_wires[16][4] ),
    .X(_01997_));
 sky130_fd_sc_hd__or2_2 _20193_ (.A(_10030_),
    .B(_11696_),
    .X(_01998_));
 sky130_fd_sc_hd__o211a_1 _20194_ (.A1(_01997_),
    .A2(_10033_),
    .B1(_01998_),
    .C1(_01840_),
    .X(_00762_));
 sky130_fd_sc_hd__buf_4 _20195_ (.A(\top_inst.grid_inst.data_path_wires[16][5] ),
    .X(_01999_));
 sky130_fd_sc_hd__or2_2 _20196_ (.A(_04858_),
    .B(_11700_),
    .X(_02000_));
 sky130_fd_sc_hd__o211a_1 _20197_ (.A1(_01999_),
    .A2(_10033_),
    .B1(_02000_),
    .C1(_01840_),
    .X(_00763_));
 sky130_fd_sc_hd__buf_4 _20198_ (.A(\top_inst.grid_inst.data_path_wires[16][6] ),
    .X(_02001_));
 sky130_fd_sc_hd__or2_2 _20199_ (.A(_04858_),
    .B(_11705_),
    .X(_02002_));
 sky130_fd_sc_hd__o211a_1 _20200_ (.A1(_02001_),
    .A2(_05739_),
    .B1(_02002_),
    .C1(_01840_),
    .X(_00764_));
 sky130_fd_sc_hd__clkbuf_4 _20201_ (.A(\top_inst.grid_inst.data_path_wires[16][7] ),
    .X(_02003_));
 sky130_fd_sc_hd__buf_4 _20202_ (.A(_02003_),
    .X(_02004_));
 sky130_fd_sc_hd__or2_2 _20203_ (.A(_04858_),
    .B(_11709_),
    .X(_02005_));
 sky130_fd_sc_hd__buf_2 _20204_ (.A(_10447_),
    .X(_02006_));
 sky130_fd_sc_hd__o211a_1 _20205_ (.A1(_02004_),
    .A2(_05739_),
    .B1(_02005_),
    .C1(_02006_),
    .X(_00765_));
 sky130_fd_sc_hd__clkbuf_4 _20206_ (.A(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[0] ),
    .X(_02007_));
 sky130_fd_sc_hd__or2_1 _20207_ (.A(_02007_),
    .B(_11689_),
    .X(_02008_));
 sky130_fd_sc_hd__o211a_1 _20208_ (.A1(_01987_),
    .A2(_11163_),
    .B1(_02008_),
    .C1(_02006_),
    .X(_00766_));
 sky130_fd_sc_hd__clkbuf_4 _20209_ (.A(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[1] ),
    .X(_02009_));
 sky130_fd_sc_hd__or2_1 _20210_ (.A(_02009_),
    .B(_11689_),
    .X(_02010_));
 sky130_fd_sc_hd__o211a_1 _20211_ (.A1(_01990_),
    .A2(_11163_),
    .B1(_02010_),
    .C1(_02006_),
    .X(_00767_));
 sky130_fd_sc_hd__clkbuf_4 _20212_ (.A(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[2] ),
    .X(_02011_));
 sky130_fd_sc_hd__or2_1 _20213_ (.A(_02011_),
    .B(_11689_),
    .X(_02012_));
 sky130_fd_sc_hd__o211a_1 _20214_ (.A1(_01993_),
    .A2(_11163_),
    .B1(_02012_),
    .C1(_02006_),
    .X(_00768_));
 sky130_fd_sc_hd__buf_4 _20215_ (.A(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[3] ),
    .X(_02013_));
 sky130_fd_sc_hd__or2_1 _20216_ (.A(_02013_),
    .B(_11689_),
    .X(_02014_));
 sky130_fd_sc_hd__o211a_1 _20217_ (.A1(_01995_),
    .A2(_11163_),
    .B1(_02014_),
    .C1(_02006_),
    .X(_00769_));
 sky130_fd_sc_hd__buf_2 _20218_ (.A(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[4] ),
    .X(_02015_));
 sky130_fd_sc_hd__clkbuf_4 _20219_ (.A(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__or2_1 _20220_ (.A(_02016_),
    .B(_11689_),
    .X(_02017_));
 sky130_fd_sc_hd__o211a_1 _20221_ (.A1(_01997_),
    .A2(_11163_),
    .B1(_02017_),
    .C1(_02006_),
    .X(_00770_));
 sky130_fd_sc_hd__clkbuf_4 _20222_ (.A(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[5] ),
    .X(_02018_));
 sky130_fd_sc_hd__or2_1 _20223_ (.A(_02018_),
    .B(_11689_),
    .X(_02019_));
 sky130_fd_sc_hd__o211a_1 _20224_ (.A1(_01999_),
    .A2(_11163_),
    .B1(_02019_),
    .C1(_02006_),
    .X(_00771_));
 sky130_fd_sc_hd__clkbuf_4 _20225_ (.A(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[6] ),
    .X(_02020_));
 sky130_fd_sc_hd__clkbuf_4 _20226_ (.A(_05772_),
    .X(_02021_));
 sky130_fd_sc_hd__or2_1 _20227_ (.A(_02020_),
    .B(_02021_),
    .X(_02022_));
 sky130_fd_sc_hd__o211a_1 _20228_ (.A1(_02001_),
    .A2(_11163_),
    .B1(_02022_),
    .C1(_02006_),
    .X(_00772_));
 sky130_fd_sc_hd__or2_1 _20229_ (.A(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[7] ),
    .B(_02021_),
    .X(_02023_));
 sky130_fd_sc_hd__o211a_1 _20230_ (.A1(_02004_),
    .A2(_11163_),
    .B1(_02023_),
    .C1(_02006_),
    .X(_00773_));
 sky130_fd_sc_hd__and3_1 _20231_ (.A(_01987_),
    .B(_02007_),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[0] ),
    .X(_02024_));
 sky130_fd_sc_hd__a21oi_1 _20232_ (.A1(_01987_),
    .A2(_02007_),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[0] ),
    .Y(_02025_));
 sky130_fd_sc_hd__o21ai_1 _20233_ (.A1(_02024_),
    .A2(_02025_),
    .B1(_08181_),
    .Y(_02026_));
 sky130_fd_sc_hd__o211a_1 _20234_ (.A1(net737),
    .A2(_01735_),
    .B1(_02026_),
    .C1(_02006_),
    .X(_00774_));
 sky130_fd_sc_hd__a22o_1 _20235_ (.A1(_01987_),
    .A2(_02009_),
    .B1(_02007_),
    .B2(_01990_),
    .X(_02027_));
 sky130_fd_sc_hd__and3_1 _20236_ (.A(_01990_),
    .B(_01987_),
    .C(_02009_),
    .X(_02028_));
 sky130_fd_sc_hd__nand2_1 _20237_ (.A(_02007_),
    .B(_02028_),
    .Y(_02029_));
 sky130_fd_sc_hd__nand3_2 _20238_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[1] ),
    .B(_02027_),
    .C(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__a21o_1 _20239_ (.A1(_02027_),
    .A2(_02029_),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[1] ),
    .X(_02031_));
 sky130_fd_sc_hd__a21oi_1 _20240_ (.A1(_02030_),
    .A2(_02031_),
    .B1(_02024_),
    .Y(_02032_));
 sky130_fd_sc_hd__and3_1 _20241_ (.A(_02024_),
    .B(_02030_),
    .C(_02031_),
    .X(_02033_));
 sky130_fd_sc_hd__o21ai_1 _20242_ (.A1(_02032_),
    .A2(_02033_),
    .B1(_06178_),
    .Y(_02034_));
 sky130_fd_sc_hd__clkbuf_4 _20243_ (.A(_10447_),
    .X(_02035_));
 sky130_fd_sc_hd__o211a_1 _20244_ (.A1(net760),
    .A2(_01735_),
    .B1(_02034_),
    .C1(_02035_),
    .X(_00775_));
 sky130_fd_sc_hd__inv_2 _20245_ (.A(_02033_),
    .Y(_02036_));
 sky130_fd_sc_hd__a22o_1 _20246_ (.A1(_01986_),
    .A2(_02011_),
    .B1(_02009_),
    .B2(_01989_),
    .X(_02037_));
 sky130_fd_sc_hd__nand4_2 _20247_ (.A(_01989_),
    .B(_01986_),
    .C(_02011_),
    .D(_02009_),
    .Y(_02038_));
 sky130_fd_sc_hd__and2_1 _20248_ (.A(_01993_),
    .B(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[0] ),
    .X(_02039_));
 sky130_fd_sc_hd__a21oi_1 _20249_ (.A1(_02037_),
    .A2(_02038_),
    .B1(_02039_),
    .Y(_02040_));
 sky130_fd_sc_hd__and3_1 _20250_ (.A(_02037_),
    .B(_02038_),
    .C(_02039_),
    .X(_02041_));
 sky130_fd_sc_hd__nor2_1 _20251_ (.A(_02040_),
    .B(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__xor2_1 _20252_ (.A(_02029_),
    .B(_02042_),
    .X(_02043_));
 sky130_fd_sc_hd__nor2_1 _20253_ (.A(_10083_),
    .B(_02043_),
    .Y(_02044_));
 sky130_fd_sc_hd__nand2_1 _20254_ (.A(_10083_),
    .B(_02043_),
    .Y(_02045_));
 sky130_fd_sc_hd__and2b_1 _20255_ (.A_N(_02044_),
    .B(_02045_),
    .X(_02046_));
 sky130_fd_sc_hd__a21oi_1 _20256_ (.A1(_02030_),
    .A2(_02036_),
    .B1(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__a31o_1 _20257_ (.A1(_02030_),
    .A2(_02036_),
    .A3(_02046_),
    .B1(_01984_),
    .X(_02048_));
 sky130_fd_sc_hd__o221a_1 _20258_ (.A1(net779),
    .A2(_01202_),
    .B1(_02047_),
    .B2(_02048_),
    .C1(_01863_),
    .X(_00776_));
 sky130_fd_sc_hd__nand2_1 _20259_ (.A(_02033_),
    .B(_02046_),
    .Y(_02049_));
 sky130_fd_sc_hd__or3b_1 _20260_ (.A(_02030_),
    .B(_02044_),
    .C_N(_02045_),
    .X(_02050_));
 sky130_fd_sc_hd__clkbuf_4 _20261_ (.A(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[2] ),
    .X(_02051_));
 sky130_fd_sc_hd__nand4_1 _20262_ (.A(_01989_),
    .B(_01986_),
    .C(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[3] ),
    .D(_02051_),
    .Y(_02052_));
 sky130_fd_sc_hd__a22o_1 _20263_ (.A1(\top_inst.grid_inst.data_path_wires[16][0] ),
    .A2(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[3] ),
    .B1(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[2] ),
    .B2(\top_inst.grid_inst.data_path_wires[16][1] ),
    .X(_02053_));
 sky130_fd_sc_hd__and4_1 _20264_ (.A(_01992_),
    .B(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[1] ),
    .C(_02052_),
    .D(_02053_),
    .X(_02054_));
 sky130_fd_sc_hd__a22o_1 _20265_ (.A1(_01992_),
    .A2(_02009_),
    .B1(_02052_),
    .B2(_02053_),
    .X(_02055_));
 sky130_fd_sc_hd__or3b_2 _20266_ (.A(_02038_),
    .B(_02054_),
    .C_N(_02055_),
    .X(_02056_));
 sky130_fd_sc_hd__nand4_1 _20267_ (.A(_01993_),
    .B(_02009_),
    .C(_02052_),
    .D(_02053_),
    .Y(_02057_));
 sky130_fd_sc_hd__a21bo_1 _20268_ (.A1(_02057_),
    .A2(_02055_),
    .B1_N(_02038_),
    .X(_02058_));
 sky130_fd_sc_hd__nand4_2 _20269_ (.A(_01995_),
    .B(_02007_),
    .C(_02056_),
    .D(_02058_),
    .Y(_02059_));
 sky130_fd_sc_hd__a22o_1 _20270_ (.A1(_01995_),
    .A2(_02007_),
    .B1(_02056_),
    .B2(_02058_),
    .X(_02060_));
 sky130_fd_sc_hd__a21oi_1 _20271_ (.A1(_02059_),
    .A2(_02060_),
    .B1(_02041_),
    .Y(_02061_));
 sky130_fd_sc_hd__and3_1 _20272_ (.A(_02041_),
    .B(_02059_),
    .C(_02060_),
    .X(_02062_));
 sky130_fd_sc_hd__or3b_1 _20273_ (.A(_02061_),
    .B(_02062_),
    .C_N(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[3] ),
    .X(_02063_));
 sky130_fd_sc_hd__o21bai_1 _20274_ (.A1(_02061_),
    .A2(_02062_),
    .B1_N(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[3] ),
    .Y(_02064_));
 sky130_fd_sc_hd__a31o_1 _20275_ (.A1(_02007_),
    .A2(_02028_),
    .A3(_02042_),
    .B1(_02044_),
    .X(_02065_));
 sky130_fd_sc_hd__and3_2 _20276_ (.A(_02063_),
    .B(_02064_),
    .C(_02065_),
    .X(_02066_));
 sky130_fd_sc_hd__a21oi_1 _20277_ (.A1(_02063_),
    .A2(_02064_),
    .B1(_02065_),
    .Y(_02067_));
 sky130_fd_sc_hd__or3_4 _20278_ (.A(_02050_),
    .B(_02066_),
    .C(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__o21ai_1 _20279_ (.A1(_02066_),
    .A2(_02067_),
    .B1(_02050_),
    .Y(_02069_));
 sky130_fd_sc_hd__nand3b_2 _20280_ (.A_N(_02049_),
    .B(_02068_),
    .C(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__a21bo_1 _20281_ (.A1(_02068_),
    .A2(_02069_),
    .B1_N(_02049_),
    .X(_02071_));
 sky130_fd_sc_hd__and2_1 _20282_ (.A(\top_inst.deskew_buff_inst.col_input[35] ),
    .B(_05730_),
    .X(_02072_));
 sky130_fd_sc_hd__a31o_1 _20283_ (.A1(_05312_),
    .A2(_02070_),
    .A3(_02071_),
    .B1(_02072_),
    .X(_02073_));
 sky130_fd_sc_hd__and2_1 _20284_ (.A(_11722_),
    .B(_02073_),
    .X(_02074_));
 sky130_fd_sc_hd__clkbuf_1 _20285_ (.A(_02074_),
    .X(_00777_));
 sky130_fd_sc_hd__and2_1 _20286_ (.A(net497),
    .B(_05634_),
    .X(_02075_));
 sky130_fd_sc_hd__nand2_2 _20287_ (.A(_01997_),
    .B(_02007_),
    .Y(_02076_));
 sky130_fd_sc_hd__and4_1 _20288_ (.A(_01989_),
    .B(_01986_),
    .C(_02013_),
    .D(_02011_),
    .X(_02077_));
 sky130_fd_sc_hd__and2_1 _20289_ (.A(\top_inst.grid_inst.data_path_wires[16][3] ),
    .B(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[1] ),
    .X(_02078_));
 sky130_fd_sc_hd__nand4_1 _20290_ (.A(_01992_),
    .B(_01989_),
    .C(_02013_),
    .D(_02011_),
    .Y(_02079_));
 sky130_fd_sc_hd__a22o_1 _20291_ (.A1(_01989_),
    .A2(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[3] ),
    .B1(_02051_),
    .B2(_01992_),
    .X(_02080_));
 sky130_fd_sc_hd__nand3_1 _20292_ (.A(_02078_),
    .B(_02079_),
    .C(_02080_),
    .Y(_02081_));
 sky130_fd_sc_hd__a21o_1 _20293_ (.A1(_02079_),
    .A2(_02080_),
    .B1(_02078_),
    .X(_02082_));
 sky130_fd_sc_hd__o211a_1 _20294_ (.A1(_02077_),
    .A2(_02054_),
    .B1(_02081_),
    .C1(_02082_),
    .X(_02083_));
 sky130_fd_sc_hd__a211o_1 _20295_ (.A1(_02081_),
    .A2(_02082_),
    .B1(_02077_),
    .C1(_02054_),
    .X(_02084_));
 sky130_fd_sc_hd__and2b_1 _20296_ (.A_N(_02083_),
    .B(_02084_),
    .X(_02085_));
 sky130_fd_sc_hd__xnor2_4 _20297_ (.A(_02076_),
    .B(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hd__nand2_2 _20298_ (.A(_02056_),
    .B(_02059_),
    .Y(_02087_));
 sky130_fd_sc_hd__xor2_4 _20299_ (.A(_02086_),
    .B(_02087_),
    .X(_02088_));
 sky130_fd_sc_hd__and3_1 _20300_ (.A(_01987_),
    .B(_02016_),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[4] ),
    .X(_02089_));
 sky130_fd_sc_hd__a21oi_1 _20301_ (.A1(_01987_),
    .A2(_02016_),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[4] ),
    .Y(_02090_));
 sky130_fd_sc_hd__or2_2 _20302_ (.A(_02089_),
    .B(_02090_),
    .X(_02091_));
 sky130_fd_sc_hd__xnor2_4 _20303_ (.A(_02088_),
    .B(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__nor2b_2 _20304_ (.A(_02062_),
    .B_N(_02063_),
    .Y(_02093_));
 sky130_fd_sc_hd__xor2_4 _20305_ (.A(_02092_),
    .B(_02093_),
    .X(_02094_));
 sky130_fd_sc_hd__o21ba_1 _20306_ (.A1(_02050_),
    .A2(_02067_),
    .B1_N(_02066_),
    .X(_02095_));
 sky130_fd_sc_hd__xnor2_2 _20307_ (.A(_02094_),
    .B(_02095_),
    .Y(_02096_));
 sky130_fd_sc_hd__a21oi_1 _20308_ (.A1(_02070_),
    .A2(_02096_),
    .B1(_05406_),
    .Y(_02097_));
 sky130_fd_sc_hd__o21a_1 _20309_ (.A1(_02070_),
    .A2(_02096_),
    .B1(_02097_),
    .X(_02098_));
 sky130_fd_sc_hd__o21a_1 _20310_ (.A1(_02075_),
    .A2(_02098_),
    .B1(_04870_),
    .X(_00778_));
 sky130_fd_sc_hd__o22ai_4 _20311_ (.A1(_02068_),
    .A2(_02094_),
    .B1(_02096_),
    .B2(_02070_),
    .Y(_02099_));
 sky130_fd_sc_hd__nand2_1 _20312_ (.A(_02086_),
    .B(_02087_),
    .Y(_02100_));
 sky130_fd_sc_hd__or3b_1 _20313_ (.A(_02089_),
    .B(_02090_),
    .C_N(_02088_),
    .X(_02101_));
 sky130_fd_sc_hd__nand3_2 _20314_ (.A(_01990_),
    .B(_02016_),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[5] ),
    .Y(_02102_));
 sky130_fd_sc_hd__a21o_1 _20315_ (.A1(_01990_),
    .A2(_02016_),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[5] ),
    .X(_02103_));
 sky130_fd_sc_hd__and3_1 _20316_ (.A(_02089_),
    .B(_02102_),
    .C(_02103_),
    .X(_02104_));
 sky130_fd_sc_hd__a21oi_1 _20317_ (.A1(_02102_),
    .A2(_02103_),
    .B1(_02089_),
    .Y(_02105_));
 sky130_fd_sc_hd__a22oi_1 _20318_ (.A1(_01987_),
    .A2(_02018_),
    .B1(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[0] ),
    .B2(_01999_),
    .Y(_02106_));
 sky130_fd_sc_hd__and4_1 _20319_ (.A(\top_inst.grid_inst.data_path_wires[16][5] ),
    .B(_01986_),
    .C(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[5] ),
    .D(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[0] ),
    .X(_02107_));
 sky130_fd_sc_hd__nor2_1 _20320_ (.A(_02106_),
    .B(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__and2_1 _20321_ (.A(\top_inst.grid_inst.data_path_wires[16][4] ),
    .B(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[1] ),
    .X(_02109_));
 sky130_fd_sc_hd__a22o_1 _20322_ (.A1(\top_inst.grid_inst.data_path_wires[16][2] ),
    .A2(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[3] ),
    .B1(_02051_),
    .B2(\top_inst.grid_inst.data_path_wires[16][3] ),
    .X(_02110_));
 sky130_fd_sc_hd__nand4_1 _20323_ (.A(\top_inst.grid_inst.data_path_wires[16][3] ),
    .B(_01992_),
    .C(_02013_),
    .D(_02051_),
    .Y(_02111_));
 sky130_fd_sc_hd__nand3_1 _20324_ (.A(_02109_),
    .B(_02110_),
    .C(_02111_),
    .Y(_02112_));
 sky130_fd_sc_hd__a21o_1 _20325_ (.A1(_02110_),
    .A2(_02111_),
    .B1(_02109_),
    .X(_02113_));
 sky130_fd_sc_hd__a21bo_1 _20326_ (.A1(_02078_),
    .A2(_02080_),
    .B1_N(_02079_),
    .X(_02114_));
 sky130_fd_sc_hd__nand3_1 _20327_ (.A(_02112_),
    .B(_02113_),
    .C(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__a21o_1 _20328_ (.A1(_02112_),
    .A2(_02113_),
    .B1(_02114_),
    .X(_02116_));
 sky130_fd_sc_hd__nand3_1 _20329_ (.A(_02108_),
    .B(_02115_),
    .C(_02116_),
    .Y(_02117_));
 sky130_fd_sc_hd__a21o_1 _20330_ (.A1(_02115_),
    .A2(_02116_),
    .B1(_02108_),
    .X(_02118_));
 sky130_fd_sc_hd__a31o_1 _20331_ (.A1(_01997_),
    .A2(_02007_),
    .A3(_02084_),
    .B1(_02083_),
    .X(_02119_));
 sky130_fd_sc_hd__nand3_2 _20332_ (.A(_02117_),
    .B(_02118_),
    .C(_02119_),
    .Y(_02120_));
 sky130_fd_sc_hd__a21o_1 _20333_ (.A1(_02117_),
    .A2(_02118_),
    .B1(_02119_),
    .X(_02121_));
 sky130_fd_sc_hd__or4bb_4 _20334_ (.A(_02104_),
    .B(_02105_),
    .C_N(_02120_),
    .D_N(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__a2bb2o_1 _20335_ (.A1_N(_02104_),
    .A2_N(_02105_),
    .B1(_02120_),
    .B2(_02121_),
    .X(_02123_));
 sky130_fd_sc_hd__nand2_1 _20336_ (.A(_02122_),
    .B(_02123_),
    .Y(_02124_));
 sky130_fd_sc_hd__a21o_1 _20337_ (.A1(_02100_),
    .A2(_02101_),
    .B1(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__nand3_1 _20338_ (.A(_02100_),
    .B(_02101_),
    .C(_02124_),
    .Y(_02126_));
 sky130_fd_sc_hd__and2_2 _20339_ (.A(_02125_),
    .B(_02126_),
    .X(_02127_));
 sky130_fd_sc_hd__xnor2_2 _20340_ (.A(_02092_),
    .B(_02093_),
    .Y(_02128_));
 sky130_fd_sc_hd__and2b_1 _20341_ (.A_N(_02093_),
    .B(_02092_),
    .X(_02129_));
 sky130_fd_sc_hd__a21oi_1 _20342_ (.A1(_02066_),
    .A2(_02128_),
    .B1(_02129_),
    .Y(_02130_));
 sky130_fd_sc_hd__xnor2_2 _20343_ (.A(_02127_),
    .B(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hd__and2_1 _20344_ (.A(_02099_),
    .B(_02131_),
    .X(_02132_));
 sky130_fd_sc_hd__o21ai_1 _20345_ (.A1(_02099_),
    .A2(_02131_),
    .B1(_05335_),
    .Y(_02133_));
 sky130_fd_sc_hd__o2bb2a_1 _20346_ (.A1_N(\top_inst.deskew_buff_inst.col_input[37] ),
    .A2_N(_05634_),
    .B1(_02132_),
    .B2(_02133_),
    .X(_02134_));
 sky130_fd_sc_hd__nor2_1 _20347_ (.A(_05440_),
    .B(_02134_),
    .Y(_00779_));
 sky130_fd_sc_hd__clkbuf_4 _20348_ (.A(_04873_),
    .X(_02135_));
 sky130_fd_sc_hd__a32oi_4 _20349_ (.A1(_02066_),
    .A2(_02128_),
    .A3(_02127_),
    .B1(_02131_),
    .B2(_02099_),
    .Y(_02136_));
 sky130_fd_sc_hd__nand3_1 _20350_ (.A(_01993_),
    .B(_02015_),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[6] ),
    .Y(_02137_));
 sky130_fd_sc_hd__a21o_1 _20351_ (.A1(_01992_),
    .A2(_02015_),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[6] ),
    .X(_02138_));
 sky130_fd_sc_hd__and3_1 _20352_ (.A(_02107_),
    .B(_02137_),
    .C(_02138_),
    .X(_02139_));
 sky130_fd_sc_hd__a21oi_1 _20353_ (.A1(_02137_),
    .A2(_02138_),
    .B1(_02107_),
    .Y(_02140_));
 sky130_fd_sc_hd__o21a_1 _20354_ (.A1(_02139_),
    .A2(_02140_),
    .B1(_02102_),
    .X(_02141_));
 sky130_fd_sc_hd__nor3_1 _20355_ (.A(_02102_),
    .B(_02139_),
    .C(_02140_),
    .Y(_02142_));
 sky130_fd_sc_hd__or2_1 _20356_ (.A(_02141_),
    .B(_02142_),
    .X(_02143_));
 sky130_fd_sc_hd__nand2_1 _20357_ (.A(_01989_),
    .B(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[5] ),
    .Y(_02144_));
 sky130_fd_sc_hd__a22oi_1 _20358_ (.A1(_01986_),
    .A2(_02020_),
    .B1(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[0] ),
    .B2(\top_inst.grid_inst.data_path_wires[16][6] ),
    .Y(_02145_));
 sky130_fd_sc_hd__and4_1 _20359_ (.A(\top_inst.grid_inst.data_path_wires[16][6] ),
    .B(_01986_),
    .C(_02020_),
    .D(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[0] ),
    .X(_02146_));
 sky130_fd_sc_hd__nor2_1 _20360_ (.A(_02145_),
    .B(_02146_),
    .Y(_02147_));
 sky130_fd_sc_hd__xnor2_1 _20361_ (.A(_02144_),
    .B(_02147_),
    .Y(_02148_));
 sky130_fd_sc_hd__and2_1 _20362_ (.A(\top_inst.grid_inst.data_path_wires[16][5] ),
    .B(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[1] ),
    .X(_02149_));
 sky130_fd_sc_hd__a22o_1 _20363_ (.A1(\top_inst.grid_inst.data_path_wires[16][3] ),
    .A2(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[3] ),
    .B1(_02051_),
    .B2(\top_inst.grid_inst.data_path_wires[16][4] ),
    .X(_02150_));
 sky130_fd_sc_hd__nand4_2 _20364_ (.A(\top_inst.grid_inst.data_path_wires[16][4] ),
    .B(\top_inst.grid_inst.data_path_wires[16][3] ),
    .C(_02013_),
    .D(_02051_),
    .Y(_02151_));
 sky130_fd_sc_hd__nand3_1 _20365_ (.A(_02149_),
    .B(_02150_),
    .C(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__a21o_1 _20366_ (.A1(_02150_),
    .A2(_02151_),
    .B1(_02149_),
    .X(_02153_));
 sky130_fd_sc_hd__a21bo_1 _20367_ (.A1(_02109_),
    .A2(_02110_),
    .B1_N(_02111_),
    .X(_02154_));
 sky130_fd_sc_hd__nand3_1 _20368_ (.A(_02152_),
    .B(_02153_),
    .C(_02154_),
    .Y(_02155_));
 sky130_fd_sc_hd__a21o_1 _20369_ (.A1(_02152_),
    .A2(_02153_),
    .B1(_02154_),
    .X(_02156_));
 sky130_fd_sc_hd__nand3_1 _20370_ (.A(_02148_),
    .B(_02155_),
    .C(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__a21o_1 _20371_ (.A1(_02155_),
    .A2(_02156_),
    .B1(_02148_),
    .X(_02158_));
 sky130_fd_sc_hd__a21bo_1 _20372_ (.A1(_02108_),
    .A2(_02116_),
    .B1_N(_02115_),
    .X(_02159_));
 sky130_fd_sc_hd__and3_1 _20373_ (.A(_02157_),
    .B(_02158_),
    .C(_02159_),
    .X(_02160_));
 sky130_fd_sc_hd__a21oi_1 _20374_ (.A1(_02157_),
    .A2(_02158_),
    .B1(_02159_),
    .Y(_02161_));
 sky130_fd_sc_hd__nor3_2 _20375_ (.A(_02143_),
    .B(_02160_),
    .C(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hd__o21a_1 _20376_ (.A1(_02160_),
    .A2(_02161_),
    .B1(_02143_),
    .X(_02163_));
 sky130_fd_sc_hd__a211oi_4 _20377_ (.A1(_02120_),
    .A2(_02122_),
    .B1(_02162_),
    .C1(_02163_),
    .Y(_02164_));
 sky130_fd_sc_hd__o211a_1 _20378_ (.A1(_02162_),
    .A2(_02163_),
    .B1(_02120_),
    .C1(_02122_),
    .X(_02165_));
 sky130_fd_sc_hd__nor3b_1 _20379_ (.A(_02164_),
    .B(_02165_),
    .C_N(_02104_),
    .Y(_02166_));
 sky130_fd_sc_hd__o21ba_1 _20380_ (.A1(_02164_),
    .A2(_02165_),
    .B1_N(_02104_),
    .X(_02167_));
 sky130_fd_sc_hd__or2_2 _20381_ (.A(_02166_),
    .B(_02167_),
    .X(_02168_));
 sky130_fd_sc_hd__a21bo_1 _20382_ (.A1(_02129_),
    .A2(_02127_),
    .B1_N(_02125_),
    .X(_02169_));
 sky130_fd_sc_hd__xor2_1 _20383_ (.A(_02168_),
    .B(_02169_),
    .X(_02170_));
 sky130_fd_sc_hd__or2_1 _20384_ (.A(_02136_),
    .B(_02170_),
    .X(_02171_));
 sky130_fd_sc_hd__a21oi_1 _20385_ (.A1(_02136_),
    .A2(_02170_),
    .B1(_05399_),
    .Y(_02172_));
 sky130_fd_sc_hd__a22o_1 _20386_ (.A1(\top_inst.deskew_buff_inst.col_input[38] ),
    .A2(_11723_),
    .B1(_02171_),
    .B2(_02172_),
    .X(_02173_));
 sky130_fd_sc_hd__and2_1 _20387_ (.A(_02135_),
    .B(_02173_),
    .X(_02174_));
 sky130_fd_sc_hd__clkbuf_1 _20388_ (.A(_02174_),
    .X(_00780_));
 sky130_fd_sc_hd__nand2_1 _20389_ (.A(_02129_),
    .B(_02127_),
    .Y(_02175_));
 sky130_fd_sc_hd__o21a_1 _20390_ (.A1(_02168_),
    .A2(_02175_),
    .B1(_02171_),
    .X(_02176_));
 sky130_fd_sc_hd__o21ba_1 _20391_ (.A1(_02144_),
    .A2(_02145_),
    .B1_N(_02146_),
    .X(_02177_));
 sky130_fd_sc_hd__inv_2 _20392_ (.A(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[7] ),
    .Y(_02178_));
 sky130_fd_sc_hd__a21oi_1 _20393_ (.A1(\top_inst.grid_inst.data_path_wires[16][3] ),
    .A2(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[7] ),
    .Y(_02179_));
 sky130_fd_sc_hd__and3_1 _20394_ (.A(\top_inst.grid_inst.data_path_wires[16][3] ),
    .B(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[4] ),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[7] ),
    .X(_02180_));
 sky130_fd_sc_hd__o22a_1 _20395_ (.A1(_01986_),
    .A2(_02178_),
    .B1(_02179_),
    .B2(_02180_),
    .X(_02181_));
 sky130_fd_sc_hd__nor4_1 _20396_ (.A(_01986_),
    .B(_02178_),
    .C(_02179_),
    .D(_02180_),
    .Y(_02182_));
 sky130_fd_sc_hd__nor2_1 _20397_ (.A(_02181_),
    .B(_02182_),
    .Y(_02183_));
 sky130_fd_sc_hd__xnor2_1 _20398_ (.A(_02177_),
    .B(_02183_),
    .Y(_02184_));
 sky130_fd_sc_hd__xor2_1 _20399_ (.A(_02137_),
    .B(_02184_),
    .X(_02185_));
 sky130_fd_sc_hd__nand2_2 _20400_ (.A(\top_inst.grid_inst.data_path_wires[16][7] ),
    .B(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[0] ),
    .Y(_02186_));
 sky130_fd_sc_hd__nand2_1 _20401_ (.A(_01989_),
    .B(_02020_),
    .Y(_02187_));
 sky130_fd_sc_hd__and3_2 _20402_ (.A(\top_inst.grid_inst.data_path_wires[16][7] ),
    .B(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[6] ),
    .C(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[0] ),
    .X(_02188_));
 sky130_fd_sc_hd__a22o_1 _20403_ (.A1(_02186_),
    .A2(_02187_),
    .B1(_02188_),
    .B2(_01989_),
    .X(_02189_));
 sky130_fd_sc_hd__nand2_1 _20404_ (.A(_01992_),
    .B(_02018_),
    .Y(_02190_));
 sky130_fd_sc_hd__xor2_2 _20405_ (.A(_02189_),
    .B(_02190_),
    .X(_02191_));
 sky130_fd_sc_hd__a22o_1 _20406_ (.A1(\top_inst.grid_inst.data_path_wires[16][4] ),
    .A2(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[3] ),
    .B1(_02051_),
    .B2(\top_inst.grid_inst.data_path_wires[16][5] ),
    .X(_02192_));
 sky130_fd_sc_hd__nand4_4 _20407_ (.A(\top_inst.grid_inst.data_path_wires[16][5] ),
    .B(\top_inst.grid_inst.data_path_wires[16][4] ),
    .C(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[3] ),
    .D(_02051_),
    .Y(_02193_));
 sky130_fd_sc_hd__nand4_2 _20408_ (.A(\top_inst.grid_inst.data_path_wires[16][6] ),
    .B(_02009_),
    .C(_02192_),
    .D(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__a22o_1 _20409_ (.A1(\top_inst.grid_inst.data_path_wires[16][6] ),
    .A2(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[1] ),
    .B1(_02192_),
    .B2(_02193_),
    .X(_02195_));
 sky130_fd_sc_hd__a21bo_1 _20410_ (.A1(_02149_),
    .A2(_02150_),
    .B1_N(_02151_),
    .X(_02196_));
 sky130_fd_sc_hd__nand3_1 _20411_ (.A(_02194_),
    .B(_02195_),
    .C(_02196_),
    .Y(_02197_));
 sky130_fd_sc_hd__a21o_1 _20412_ (.A1(_02194_),
    .A2(_02195_),
    .B1(_02196_),
    .X(_02198_));
 sky130_fd_sc_hd__nand3_1 _20413_ (.A(_02191_),
    .B(_02197_),
    .C(_02198_),
    .Y(_02199_));
 sky130_fd_sc_hd__a21o_1 _20414_ (.A1(_02197_),
    .A2(_02198_),
    .B1(_02191_),
    .X(_02200_));
 sky130_fd_sc_hd__a21bo_1 _20415_ (.A1(_02148_),
    .A2(_02156_),
    .B1_N(_02155_),
    .X(_02201_));
 sky130_fd_sc_hd__and3_1 _20416_ (.A(_02199_),
    .B(_02200_),
    .C(_02201_),
    .X(_02202_));
 sky130_fd_sc_hd__a21oi_1 _20417_ (.A1(_02199_),
    .A2(_02200_),
    .B1(_02201_),
    .Y(_02203_));
 sky130_fd_sc_hd__or3_1 _20418_ (.A(_02185_),
    .B(_02202_),
    .C(_02203_),
    .X(_02204_));
 sky130_fd_sc_hd__o21ai_1 _20419_ (.A1(_02202_),
    .A2(_02203_),
    .B1(_02185_),
    .Y(_02205_));
 sky130_fd_sc_hd__o211ai_2 _20420_ (.A1(_02160_),
    .A2(_02162_),
    .B1(_02204_),
    .C1(_02205_),
    .Y(_02206_));
 sky130_fd_sc_hd__a211o_1 _20421_ (.A1(_02204_),
    .A2(_02205_),
    .B1(_02160_),
    .C1(_02162_),
    .X(_02207_));
 sky130_fd_sc_hd__o211ai_2 _20422_ (.A1(_02139_),
    .A2(_02142_),
    .B1(_02206_),
    .C1(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__a211o_1 _20423_ (.A1(_02206_),
    .A2(_02207_),
    .B1(_02139_),
    .C1(_02142_),
    .X(_02209_));
 sky130_fd_sc_hd__o211ai_2 _20424_ (.A1(_02164_),
    .A2(_02166_),
    .B1(_02208_),
    .C1(_02209_),
    .Y(_02210_));
 sky130_fd_sc_hd__a211o_1 _20425_ (.A1(_02208_),
    .A2(_02209_),
    .B1(_02164_),
    .C1(_02166_),
    .X(_02211_));
 sky130_fd_sc_hd__and3_1 _20426_ (.A(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[7] ),
    .B(_02210_),
    .C(_02211_),
    .X(_02212_));
 sky130_fd_sc_hd__a21oi_1 _20427_ (.A1(_02210_),
    .A2(_02211_),
    .B1(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[7] ),
    .Y(_02213_));
 sky130_fd_sc_hd__nor2_1 _20428_ (.A(_02125_),
    .B(_02168_),
    .Y(_02214_));
 sky130_fd_sc_hd__o21ba_1 _20429_ (.A1(_02212_),
    .A2(_02213_),
    .B1_N(_02214_),
    .X(_02215_));
 sky130_fd_sc_hd__or3b_1 _20430_ (.A(_02212_),
    .B(_02213_),
    .C_N(_02214_),
    .X(_02216_));
 sky130_fd_sc_hd__or2b_1 _20431_ (.A(_02215_),
    .B_N(_02216_),
    .X(_02217_));
 sky130_fd_sc_hd__xnor2_1 _20432_ (.A(_02176_),
    .B(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__nand2_1 _20433_ (.A(_05317_),
    .B(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__o211a_1 _20434_ (.A1(net745),
    .A2(_01735_),
    .B1(_02219_),
    .C1(_02035_),
    .X(_00781_));
 sky130_fd_sc_hd__o221a_1 _20435_ (.A1(_02168_),
    .A2(_02175_),
    .B1(_02170_),
    .B2(_02136_),
    .C1(_02216_),
    .X(_02220_));
 sky130_fd_sc_hd__nor2_1 _20436_ (.A(_02215_),
    .B(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__nand2_1 _20437_ (.A(_02206_),
    .B(_02208_),
    .Y(_02222_));
 sky130_fd_sc_hd__and2b_1 _20438_ (.A_N(_02177_),
    .B(_02183_),
    .X(_02223_));
 sky130_fd_sc_hd__a41o_1 _20439_ (.A1(_01993_),
    .A2(_02016_),
    .A3(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[6] ),
    .A4(_02184_),
    .B1(_02223_),
    .X(_02224_));
 sky130_fd_sc_hd__nor3_1 _20440_ (.A(_02185_),
    .B(_02202_),
    .C(_02203_),
    .Y(_02225_));
 sky130_fd_sc_hd__nor2_1 _20441_ (.A(_02180_),
    .B(_02182_),
    .Y(_02226_));
 sky130_fd_sc_hd__clkbuf_4 _20442_ (.A(_02188_),
    .X(_02227_));
 sky130_fd_sc_hd__o2bb2a_1 _20443_ (.A1_N(_01990_),
    .A2_N(_02227_),
    .B1(_02189_),
    .B2(_02190_),
    .X(_02228_));
 sky130_fd_sc_hd__clkbuf_4 _20444_ (.A(_02178_),
    .X(_02229_));
 sky130_fd_sc_hd__a21oi_1 _20445_ (.A1(\top_inst.grid_inst.data_path_wires[16][4] ),
    .A2(_02015_),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[8] ),
    .Y(_02230_));
 sky130_fd_sc_hd__and3_1 _20446_ (.A(\top_inst.grid_inst.data_path_wires[16][4] ),
    .B(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[4] ),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[8] ),
    .X(_02231_));
 sky130_fd_sc_hd__o22a_1 _20447_ (.A1(_01990_),
    .A2(_02229_),
    .B1(_02230_),
    .B2(_02231_),
    .X(_02232_));
 sky130_fd_sc_hd__nor4_1 _20448_ (.A(_01990_),
    .B(_02229_),
    .C(_02230_),
    .D(_02231_),
    .Y(_02233_));
 sky130_fd_sc_hd__nor2_1 _20449_ (.A(_02232_),
    .B(net179),
    .Y(_02234_));
 sky130_fd_sc_hd__xnor2_1 _20450_ (.A(_02228_),
    .B(_02234_),
    .Y(_02235_));
 sky130_fd_sc_hd__xnor2_1 _20451_ (.A(_02226_),
    .B(_02235_),
    .Y(_02236_));
 sky130_fd_sc_hd__nand2_1 _20452_ (.A(_01992_),
    .B(_02020_),
    .Y(_02237_));
 sky130_fd_sc_hd__a22o_1 _20453_ (.A1(_01992_),
    .A2(_02188_),
    .B1(_02237_),
    .B2(_02186_),
    .X(_02238_));
 sky130_fd_sc_hd__nand2_1 _20454_ (.A(_01995_),
    .B(_02018_),
    .Y(_02239_));
 sky130_fd_sc_hd__xor2_2 _20455_ (.A(_02238_),
    .B(_02239_),
    .X(_02240_));
 sky130_fd_sc_hd__and2_1 _20456_ (.A(_02003_),
    .B(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[1] ),
    .X(_02241_));
 sky130_fd_sc_hd__a22o_1 _20457_ (.A1(\top_inst.grid_inst.data_path_wires[16][5] ),
    .A2(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[3] ),
    .B1(_02051_),
    .B2(\top_inst.grid_inst.data_path_wires[16][6] ),
    .X(_02242_));
 sky130_fd_sc_hd__nand4_1 _20458_ (.A(\top_inst.grid_inst.data_path_wires[16][6] ),
    .B(\top_inst.grid_inst.data_path_wires[16][5] ),
    .C(_02013_),
    .D(_02011_),
    .Y(_02243_));
 sky130_fd_sc_hd__and3_1 _20459_ (.A(_02241_),
    .B(_02242_),
    .C(_02243_),
    .X(_02244_));
 sky130_fd_sc_hd__a21oi_1 _20460_ (.A1(_02242_),
    .A2(_02243_),
    .B1(_02241_),
    .Y(_02245_));
 sky130_fd_sc_hd__a211o_1 _20461_ (.A1(_02193_),
    .A2(_02194_),
    .B1(_02244_),
    .C1(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__o211ai_2 _20462_ (.A1(_02244_),
    .A2(_02245_),
    .B1(_02193_),
    .C1(_02194_),
    .Y(_02247_));
 sky130_fd_sc_hd__nand3_1 _20463_ (.A(_02240_),
    .B(_02246_),
    .C(_02247_),
    .Y(_02248_));
 sky130_fd_sc_hd__a21o_1 _20464_ (.A1(_02246_),
    .A2(_02247_),
    .B1(_02240_),
    .X(_02249_));
 sky130_fd_sc_hd__a21bo_1 _20465_ (.A1(_02191_),
    .A2(_02198_),
    .B1_N(_02197_),
    .X(_02250_));
 sky130_fd_sc_hd__nand3_2 _20466_ (.A(_02248_),
    .B(_02249_),
    .C(_02250_),
    .Y(_02251_));
 sky130_fd_sc_hd__a21o_1 _20467_ (.A1(_02248_),
    .A2(_02249_),
    .B1(_02250_),
    .X(_02252_));
 sky130_fd_sc_hd__nand3_1 _20468_ (.A(_02236_),
    .B(_02251_),
    .C(_02252_),
    .Y(_02253_));
 sky130_fd_sc_hd__a21o_1 _20469_ (.A1(_02251_),
    .A2(_02252_),
    .B1(_02236_),
    .X(_02254_));
 sky130_fd_sc_hd__o211ai_2 _20470_ (.A1(_02202_),
    .A2(_02225_),
    .B1(_02253_),
    .C1(_02254_),
    .Y(_02255_));
 sky130_fd_sc_hd__a211o_1 _20471_ (.A1(_02253_),
    .A2(_02254_),
    .B1(_02202_),
    .C1(_02225_),
    .X(_02256_));
 sky130_fd_sc_hd__and3_1 _20472_ (.A(_02224_),
    .B(_02255_),
    .C(_02256_),
    .X(_02257_));
 sky130_fd_sc_hd__a21oi_1 _20473_ (.A1(_02255_),
    .A2(_02256_),
    .B1(_02224_),
    .Y(_02258_));
 sky130_fd_sc_hd__nor2_1 _20474_ (.A(_02257_),
    .B(_02258_),
    .Y(_02259_));
 sky130_fd_sc_hd__xnor2_1 _20475_ (.A(_02222_),
    .B(_02259_),
    .Y(_02260_));
 sky130_fd_sc_hd__a21boi_1 _20476_ (.A1(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[7] ),
    .A2(_02211_),
    .B1_N(_02210_),
    .Y(_02261_));
 sky130_fd_sc_hd__xnor2_1 _20477_ (.A(_02260_),
    .B(_02261_),
    .Y(_02262_));
 sky130_fd_sc_hd__inv_2 _20478_ (.A(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__nand2_1 _20479_ (.A(_02221_),
    .B(_02263_),
    .Y(_02264_));
 sky130_fd_sc_hd__or2_1 _20480_ (.A(_02221_),
    .B(_02263_),
    .X(_02265_));
 sky130_fd_sc_hd__a21o_1 _20481_ (.A1(_02264_),
    .A2(_02265_),
    .B1(_05732_),
    .X(_02266_));
 sky130_fd_sc_hd__o211a_1 _20482_ (.A1(net871),
    .A2(_01735_),
    .B1(_02266_),
    .C1(_02035_),
    .X(_00782_));
 sky130_fd_sc_hd__or2_1 _20483_ (.A(_02260_),
    .B(_02261_),
    .X(_02267_));
 sky130_fd_sc_hd__nand2_1 _20484_ (.A(_02267_),
    .B(_02264_),
    .Y(_02268_));
 sky130_fd_sc_hd__nand2_1 _20485_ (.A(_02222_),
    .B(_02259_),
    .Y(_02269_));
 sky130_fd_sc_hd__or2b_1 _20486_ (.A(_02226_),
    .B_N(_02235_),
    .X(_02270_));
 sky130_fd_sc_hd__o31ai_2 _20487_ (.A1(_02228_),
    .A2(_02232_),
    .A3(net178),
    .B1(_02270_),
    .Y(_02271_));
 sky130_fd_sc_hd__inv_2 _20488_ (.A(_02251_),
    .Y(_02272_));
 sky130_fd_sc_hd__and3_1 _20489_ (.A(_02236_),
    .B(_02251_),
    .C(_02252_),
    .X(_02273_));
 sky130_fd_sc_hd__or2_1 _20490_ (.A(_02231_),
    .B(_02233_),
    .X(_02274_));
 sky130_fd_sc_hd__o2bb2a_1 _20491_ (.A1_N(_01993_),
    .A2_N(_02227_),
    .B1(_02238_),
    .B2(_02239_),
    .X(_02275_));
 sky130_fd_sc_hd__a21oi_1 _20492_ (.A1(_01999_),
    .A2(_02015_),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[9] ),
    .Y(_02276_));
 sky130_fd_sc_hd__and3_1 _20493_ (.A(\top_inst.grid_inst.data_path_wires[16][5] ),
    .B(_02015_),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[9] ),
    .X(_02277_));
 sky130_fd_sc_hd__o22a_1 _20494_ (.A1(_01993_),
    .A2(_02229_),
    .B1(_02276_),
    .B2(_02277_),
    .X(_02278_));
 sky130_fd_sc_hd__nor4_1 _20495_ (.A(_01993_),
    .B(_02229_),
    .C(_02276_),
    .D(_02277_),
    .Y(_02279_));
 sky130_fd_sc_hd__nor2_1 _20496_ (.A(_02278_),
    .B(_02279_),
    .Y(_02280_));
 sky130_fd_sc_hd__xnor2_1 _20497_ (.A(_02275_),
    .B(_02280_),
    .Y(_02281_));
 sky130_fd_sc_hd__xor2_1 _20498_ (.A(_02274_),
    .B(_02281_),
    .X(_02282_));
 sky130_fd_sc_hd__nand2_1 _20499_ (.A(\top_inst.grid_inst.data_path_wires[16][3] ),
    .B(_02020_),
    .Y(_02283_));
 sky130_fd_sc_hd__a22o_1 _20500_ (.A1(_01995_),
    .A2(_02188_),
    .B1(_02283_),
    .B2(_02186_),
    .X(_02284_));
 sky130_fd_sc_hd__nand2_1 _20501_ (.A(_01997_),
    .B(_02018_),
    .Y(_02285_));
 sky130_fd_sc_hd__xor2_2 _20502_ (.A(_02284_),
    .B(_02285_),
    .X(_02286_));
 sky130_fd_sc_hd__and4_1 _20503_ (.A(\top_inst.grid_inst.data_path_wires[16][6] ),
    .B(\top_inst.grid_inst.data_path_wires[16][5] ),
    .C(_02013_),
    .D(_02011_),
    .X(_02287_));
 sky130_fd_sc_hd__a22oi_2 _20504_ (.A1(\top_inst.grid_inst.data_path_wires[16][6] ),
    .A2(_02013_),
    .B1(_02011_),
    .B2(_02003_),
    .Y(_02288_));
 sky130_fd_sc_hd__and4_1 _20505_ (.A(_02003_),
    .B(\top_inst.grid_inst.data_path_wires[16][6] ),
    .C(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[3] ),
    .D(_02051_),
    .X(_02289_));
 sky130_fd_sc_hd__o21a_1 _20506_ (.A1(_02288_),
    .A2(_02289_),
    .B1(_02241_),
    .X(_02290_));
 sky130_fd_sc_hd__nor3_1 _20507_ (.A(_02241_),
    .B(_02288_),
    .C(_02289_),
    .Y(_02291_));
 sky130_fd_sc_hd__o22ai_2 _20508_ (.A1(_02287_),
    .A2(_02244_),
    .B1(_02290_),
    .B2(_02291_),
    .Y(_02292_));
 sky130_fd_sc_hd__or4_2 _20509_ (.A(_02287_),
    .B(_02244_),
    .C(_02290_),
    .D(_02291_),
    .X(_02293_));
 sky130_fd_sc_hd__nand3_1 _20510_ (.A(_02286_),
    .B(_02292_),
    .C(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__a21o_1 _20511_ (.A1(_02292_),
    .A2(_02293_),
    .B1(_02286_),
    .X(_02295_));
 sky130_fd_sc_hd__a21bo_1 _20512_ (.A1(_02240_),
    .A2(_02247_),
    .B1_N(_02246_),
    .X(_02296_));
 sky130_fd_sc_hd__nand3_2 _20513_ (.A(_02294_),
    .B(_02295_),
    .C(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__a21o_1 _20514_ (.A1(_02294_),
    .A2(_02295_),
    .B1(_02296_),
    .X(_02298_));
 sky130_fd_sc_hd__nand3_2 _20515_ (.A(_02282_),
    .B(_02297_),
    .C(_02298_),
    .Y(_02299_));
 sky130_fd_sc_hd__a21o_1 _20516_ (.A1(_02297_),
    .A2(_02298_),
    .B1(_02282_),
    .X(_02300_));
 sky130_fd_sc_hd__o211ai_2 _20517_ (.A1(_02272_),
    .A2(_02273_),
    .B1(_02299_),
    .C1(_02300_),
    .Y(_02301_));
 sky130_fd_sc_hd__a211o_1 _20518_ (.A1(_02299_),
    .A2(_02300_),
    .B1(_02272_),
    .C1(_02273_),
    .X(_02302_));
 sky130_fd_sc_hd__and3_1 _20519_ (.A(_02271_),
    .B(_02301_),
    .C(_02302_),
    .X(_02303_));
 sky130_fd_sc_hd__a21oi_1 _20520_ (.A1(_02301_),
    .A2(_02302_),
    .B1(_02271_),
    .Y(_02304_));
 sky130_fd_sc_hd__nor2_1 _20521_ (.A(_02303_),
    .B(_02304_),
    .Y(_02305_));
 sky130_fd_sc_hd__a21bo_1 _20522_ (.A1(_02224_),
    .A2(_02256_),
    .B1_N(_02255_),
    .X(_02306_));
 sky130_fd_sc_hd__xnor2_2 _20523_ (.A(_02305_),
    .B(_02306_),
    .Y(_02307_));
 sky130_fd_sc_hd__xnor2_2 _20524_ (.A(_02269_),
    .B(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__a21oi_1 _20525_ (.A1(_02268_),
    .A2(_02308_),
    .B1(_07576_),
    .Y(_02309_));
 sky130_fd_sc_hd__o21ai_1 _20526_ (.A1(_02268_),
    .A2(_02308_),
    .B1(_02309_),
    .Y(_02310_));
 sky130_fd_sc_hd__o211a_1 _20527_ (.A1(net883),
    .A2(_01735_),
    .B1(_02310_),
    .C1(_02035_),
    .X(_00783_));
 sky130_fd_sc_hd__nand2_1 _20528_ (.A(_02305_),
    .B(_02306_),
    .Y(_02311_));
 sky130_fd_sc_hd__a21bo_1 _20529_ (.A1(_02271_),
    .A2(_02302_),
    .B1_N(_02301_),
    .X(_02312_));
 sky130_fd_sc_hd__nand2_1 _20530_ (.A(_02274_),
    .B(_02281_),
    .Y(_02313_));
 sky130_fd_sc_hd__o31ai_4 _20531_ (.A1(_02275_),
    .A2(_02278_),
    .A3(net177),
    .B1(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__or2_1 _20532_ (.A(_02277_),
    .B(_02279_),
    .X(_02315_));
 sky130_fd_sc_hd__o2bb2a_1 _20533_ (.A1_N(_01995_),
    .A2_N(_02227_),
    .B1(_02284_),
    .B2(_02285_),
    .X(_02316_));
 sky130_fd_sc_hd__a21oi_1 _20534_ (.A1(_02001_),
    .A2(_02015_),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[10] ),
    .Y(_02317_));
 sky130_fd_sc_hd__and3_1 _20535_ (.A(_02001_),
    .B(_02015_),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[10] ),
    .X(_02318_));
 sky130_fd_sc_hd__o22a_1 _20536_ (.A1(_01995_),
    .A2(_02229_),
    .B1(_02317_),
    .B2(_02318_),
    .X(_02319_));
 sky130_fd_sc_hd__nor4_1 _20537_ (.A(_01995_),
    .B(_02229_),
    .C(_02317_),
    .D(_02318_),
    .Y(_02320_));
 sky130_fd_sc_hd__nor2_1 _20538_ (.A(_02319_),
    .B(net176),
    .Y(_02321_));
 sky130_fd_sc_hd__xnor2_1 _20539_ (.A(_02316_),
    .B(_02321_),
    .Y(_02322_));
 sky130_fd_sc_hd__xor2_1 _20540_ (.A(_02315_),
    .B(_02322_),
    .X(_02323_));
 sky130_fd_sc_hd__nand2_1 _20541_ (.A(\top_inst.grid_inst.data_path_wires[16][4] ),
    .B(_02020_),
    .Y(_02324_));
 sky130_fd_sc_hd__a22o_1 _20542_ (.A1(_01997_),
    .A2(_02188_),
    .B1(_02324_),
    .B2(_02186_),
    .X(_02325_));
 sky130_fd_sc_hd__nand2_1 _20543_ (.A(_01999_),
    .B(_02018_),
    .Y(_02326_));
 sky130_fd_sc_hd__xor2_1 _20544_ (.A(_02325_),
    .B(_02326_),
    .X(_02327_));
 sky130_fd_sc_hd__o21ai_1 _20545_ (.A1(_02013_),
    .A2(_02011_),
    .B1(_02003_),
    .Y(_02328_));
 sky130_fd_sc_hd__and3_1 _20546_ (.A(_02003_),
    .B(_02013_),
    .C(_02011_),
    .X(_02329_));
 sky130_fd_sc_hd__or2_1 _20547_ (.A(_02328_),
    .B(_02329_),
    .X(_02330_));
 sky130_fd_sc_hd__inv_2 _20548_ (.A(_02009_),
    .Y(_02331_));
 sky130_fd_sc_hd__o22a_1 _20549_ (.A1(_02331_),
    .A2(_02288_),
    .B1(_02289_),
    .B2(_02241_),
    .X(_02332_));
 sky130_fd_sc_hd__xnor2_2 _20550_ (.A(_02330_),
    .B(_02332_),
    .Y(_02333_));
 sky130_fd_sc_hd__xor2_1 _20551_ (.A(_02327_),
    .B(_02333_),
    .X(_02334_));
 sky130_fd_sc_hd__a21bo_1 _20552_ (.A1(_02286_),
    .A2(_02293_),
    .B1_N(_02292_),
    .X(_02335_));
 sky130_fd_sc_hd__xor2_1 _20553_ (.A(_02334_),
    .B(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__xnor2_1 _20554_ (.A(_02323_),
    .B(_02336_),
    .Y(_02337_));
 sky130_fd_sc_hd__a21o_1 _20555_ (.A1(_02297_),
    .A2(_02299_),
    .B1(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__nand3_1 _20556_ (.A(_02297_),
    .B(_02299_),
    .C(_02337_),
    .Y(_02339_));
 sky130_fd_sc_hd__and2_1 _20557_ (.A(_02338_),
    .B(_02339_),
    .X(_02340_));
 sky130_fd_sc_hd__xor2_2 _20558_ (.A(_02314_),
    .B(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__xnor2_2 _20559_ (.A(_02312_),
    .B(_02341_),
    .Y(_02342_));
 sky130_fd_sc_hd__xor2_2 _20560_ (.A(_02311_),
    .B(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__a21o_1 _20561_ (.A1(_02269_),
    .A2(_02267_),
    .B1(_02307_),
    .X(_02344_));
 sky130_fd_sc_hd__o21ai_2 _20562_ (.A1(_02264_),
    .A2(_02308_),
    .B1(_02344_),
    .Y(_02345_));
 sky130_fd_sc_hd__nand2_1 _20563_ (.A(_02343_),
    .B(_02345_),
    .Y(_02346_));
 sky130_fd_sc_hd__o21a_1 _20564_ (.A1(_02343_),
    .A2(_02345_),
    .B1(_10831_),
    .X(_02347_));
 sky130_fd_sc_hd__a22o_1 _20565_ (.A1(\top_inst.deskew_buff_inst.col_input[42] ),
    .A2(_11723_),
    .B1(_02346_),
    .B2(_02347_),
    .X(_02348_));
 sky130_fd_sc_hd__and2_1 _20566_ (.A(_02135_),
    .B(_02348_),
    .X(_02349_));
 sky130_fd_sc_hd__clkbuf_1 _20567_ (.A(_02349_),
    .X(_00784_));
 sky130_fd_sc_hd__nor2_1 _20568_ (.A(_02311_),
    .B(_02342_),
    .Y(_02350_));
 sky130_fd_sc_hd__a21oi_1 _20569_ (.A1(_02343_),
    .A2(_02345_),
    .B1(_02350_),
    .Y(_02351_));
 sky130_fd_sc_hd__and2_1 _20570_ (.A(_02312_),
    .B(_02341_),
    .X(_02352_));
 sky130_fd_sc_hd__nand2_1 _20571_ (.A(_02315_),
    .B(_02322_),
    .Y(_02353_));
 sky130_fd_sc_hd__o31ai_2 _20572_ (.A1(_02316_),
    .A2(_02319_),
    .A3(net175),
    .B1(_02353_),
    .Y(_02354_));
 sky130_fd_sc_hd__nor2_1 _20573_ (.A(_02318_),
    .B(_02320_),
    .Y(_02355_));
 sky130_fd_sc_hd__o2bb2a_1 _20574_ (.A1_N(_01997_),
    .A2_N(_02227_),
    .B1(_02325_),
    .B2(_02326_),
    .X(_02356_));
 sky130_fd_sc_hd__a21oi_1 _20575_ (.A1(_02004_),
    .A2(_02016_),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[11] ),
    .Y(_02357_));
 sky130_fd_sc_hd__and3_1 _20576_ (.A(_02004_),
    .B(_02015_),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[11] ),
    .X(_02358_));
 sky130_fd_sc_hd__o22a_1 _20577_ (.A1(_01997_),
    .A2(_02229_),
    .B1(_02357_),
    .B2(_02358_),
    .X(_02359_));
 sky130_fd_sc_hd__nor4_1 _20578_ (.A(_01997_),
    .B(_02229_),
    .C(_02357_),
    .D(_02358_),
    .Y(_02360_));
 sky130_fd_sc_hd__nor2_1 _20579_ (.A(_02359_),
    .B(net174),
    .Y(_02361_));
 sky130_fd_sc_hd__xnor2_1 _20580_ (.A(_02356_),
    .B(_02361_),
    .Y(_02362_));
 sky130_fd_sc_hd__xnor2_1 _20581_ (.A(_02355_),
    .B(_02362_),
    .Y(_02363_));
 sky130_fd_sc_hd__and2_2 _20582_ (.A(_02009_),
    .B(_02329_),
    .X(_02364_));
 sky130_fd_sc_hd__or2b_2 _20583_ (.A(_02241_),
    .B_N(_02328_),
    .X(_02365_));
 sky130_fd_sc_hd__nand2b_2 _20584_ (.A_N(_02364_),
    .B(_02365_),
    .Y(_02366_));
 sky130_fd_sc_hd__nand2_1 _20585_ (.A(_01999_),
    .B(_02020_),
    .Y(_02367_));
 sky130_fd_sc_hd__a22o_1 _20586_ (.A1(_01999_),
    .A2(_02227_),
    .B1(_02367_),
    .B2(_02186_),
    .X(_02368_));
 sky130_fd_sc_hd__nand2_1 _20587_ (.A(_02001_),
    .B(_02018_),
    .Y(_02369_));
 sky130_fd_sc_hd__xor2_1 _20588_ (.A(_02368_),
    .B(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__xnor2_1 _20589_ (.A(_02366_),
    .B(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__a21oi_1 _20590_ (.A1(_02327_),
    .A2(_02333_),
    .B1(_02364_),
    .Y(_02372_));
 sky130_fd_sc_hd__xnor2_1 _20591_ (.A(_02371_),
    .B(_02372_),
    .Y(_02373_));
 sky130_fd_sc_hd__xnor2_1 _20592_ (.A(_02363_),
    .B(_02373_),
    .Y(_02374_));
 sky130_fd_sc_hd__and2_1 _20593_ (.A(_02334_),
    .B(_02335_),
    .X(_02375_));
 sky130_fd_sc_hd__a21o_1 _20594_ (.A1(_02323_),
    .A2(_02336_),
    .B1(_02375_),
    .X(_02376_));
 sky130_fd_sc_hd__xnor2_1 _20595_ (.A(_02374_),
    .B(_02376_),
    .Y(_02377_));
 sky130_fd_sc_hd__xnor2_1 _20596_ (.A(_02354_),
    .B(_02377_),
    .Y(_02378_));
 sky130_fd_sc_hd__a21bo_1 _20597_ (.A1(_02314_),
    .A2(_02340_),
    .B1_N(_02338_),
    .X(_02379_));
 sky130_fd_sc_hd__xnor2_1 _20598_ (.A(_02378_),
    .B(_02379_),
    .Y(_02380_));
 sky130_fd_sc_hd__xor2_1 _20599_ (.A(_02352_),
    .B(_02380_),
    .X(_02381_));
 sky130_fd_sc_hd__a21oi_1 _20600_ (.A1(_02351_),
    .A2(_02381_),
    .B1(_07576_),
    .Y(_02382_));
 sky130_fd_sc_hd__o21ai_1 _20601_ (.A1(_02351_),
    .A2(_02381_),
    .B1(_02382_),
    .Y(_02383_));
 sky130_fd_sc_hd__o211a_1 _20602_ (.A1(net795),
    .A2(_01735_),
    .B1(_02383_),
    .C1(_02035_),
    .X(_00785_));
 sky130_fd_sc_hd__nand2_1 _20603_ (.A(_02343_),
    .B(_02381_),
    .Y(_02384_));
 sky130_fd_sc_hd__or2_1 _20604_ (.A(_02344_),
    .B(_02384_),
    .X(_02385_));
 sky130_fd_sc_hd__or2_1 _20605_ (.A(_02262_),
    .B(_02308_),
    .X(_02386_));
 sky130_fd_sc_hd__o21ai_1 _20606_ (.A1(_02352_),
    .A2(_02350_),
    .B1(_02380_),
    .Y(_02387_));
 sky130_fd_sc_hd__o41a_1 _20607_ (.A1(_02215_),
    .A2(_02220_),
    .A3(_02386_),
    .A4(_02384_),
    .B1(_02387_),
    .X(_02388_));
 sky130_fd_sc_hd__nand2_1 _20608_ (.A(_02385_),
    .B(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__and2b_1 _20609_ (.A_N(_02378_),
    .B(_02379_),
    .X(_02390_));
 sky130_fd_sc_hd__or2b_1 _20610_ (.A(_02374_),
    .B_N(_02376_),
    .X(_02391_));
 sky130_fd_sc_hd__nand2_1 _20611_ (.A(_02354_),
    .B(_02377_),
    .Y(_02392_));
 sky130_fd_sc_hd__or2b_1 _20612_ (.A(_02355_),
    .B_N(_02362_),
    .X(_02393_));
 sky130_fd_sc_hd__o31a_1 _20613_ (.A1(_02356_),
    .A2(_02359_),
    .A3(net174),
    .B1(_02393_),
    .X(_02394_));
 sky130_fd_sc_hd__or2_1 _20614_ (.A(_02358_),
    .B(_02360_),
    .X(_02395_));
 sky130_fd_sc_hd__o2bb2ai_1 _20615_ (.A1_N(_01999_),
    .A2_N(_02227_),
    .B1(_02368_),
    .B2(_02369_),
    .Y(_02396_));
 sky130_fd_sc_hd__nand3_1 _20616_ (.A(_02004_),
    .B(_02016_),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[12] ),
    .Y(_02397_));
 sky130_fd_sc_hd__a21o_1 _20617_ (.A1(_02003_),
    .A2(_02015_),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[12] ),
    .X(_02398_));
 sky130_fd_sc_hd__nand2_1 _20618_ (.A(_02397_),
    .B(_02398_),
    .Y(_02399_));
 sky130_fd_sc_hd__nor2_1 _20619_ (.A(_01999_),
    .B(_02229_),
    .Y(_02400_));
 sky130_fd_sc_hd__xnor2_1 _20620_ (.A(_02399_),
    .B(_02400_),
    .Y(_02401_));
 sky130_fd_sc_hd__xor2_1 _20621_ (.A(_02396_),
    .B(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__xor2_1 _20622_ (.A(_02395_),
    .B(_02402_),
    .X(_02403_));
 sky130_fd_sc_hd__nand2_1 _20623_ (.A(_02001_),
    .B(_02020_),
    .Y(_02404_));
 sky130_fd_sc_hd__a22o_1 _20624_ (.A1(_02001_),
    .A2(_02227_),
    .B1(_02404_),
    .B2(_02186_),
    .X(_02405_));
 sky130_fd_sc_hd__nand2_2 _20625_ (.A(_02003_),
    .B(_02018_),
    .Y(_02406_));
 sky130_fd_sc_hd__xor2_1 _20626_ (.A(_02405_),
    .B(_02406_),
    .X(_02407_));
 sky130_fd_sc_hd__xnor2_1 _20627_ (.A(_02366_),
    .B(_02407_),
    .Y(_02408_));
 sky130_fd_sc_hd__a21o_1 _20628_ (.A1(_02365_),
    .A2(_02370_),
    .B1(_02364_),
    .X(_02409_));
 sky130_fd_sc_hd__xor2_1 _20629_ (.A(_02408_),
    .B(_02409_),
    .X(_02410_));
 sky130_fd_sc_hd__xnor2_1 _20630_ (.A(_02403_),
    .B(_02410_),
    .Y(_02411_));
 sky130_fd_sc_hd__and2b_1 _20631_ (.A_N(_02372_),
    .B(_02371_),
    .X(_02412_));
 sky130_fd_sc_hd__a21oi_1 _20632_ (.A1(_02363_),
    .A2(_02373_),
    .B1(_02412_),
    .Y(_02413_));
 sky130_fd_sc_hd__xnor2_1 _20633_ (.A(_02411_),
    .B(_02413_),
    .Y(_02414_));
 sky130_fd_sc_hd__xnor2_1 _20634_ (.A(_02394_),
    .B(_02414_),
    .Y(_02415_));
 sky130_fd_sc_hd__a21o_1 _20635_ (.A1(_02391_),
    .A2(_02392_),
    .B1(_02415_),
    .X(_02416_));
 sky130_fd_sc_hd__nand3_1 _20636_ (.A(_02391_),
    .B(_02392_),
    .C(_02415_),
    .Y(_02417_));
 sky130_fd_sc_hd__and2_1 _20637_ (.A(_02416_),
    .B(_02417_),
    .X(_02418_));
 sky130_fd_sc_hd__xor2_2 _20638_ (.A(_02390_),
    .B(_02418_),
    .X(_02419_));
 sky130_fd_sc_hd__xor2_1 _20639_ (.A(_02389_),
    .B(_02419_),
    .X(_02420_));
 sky130_fd_sc_hd__or2_1 _20640_ (.A(net816),
    .B(_01386_),
    .X(_02421_));
 sky130_fd_sc_hd__o211a_1 _20641_ (.A1(_01819_),
    .A2(_02420_),
    .B1(_02421_),
    .C1(_02035_),
    .X(_00786_));
 sky130_fd_sc_hd__nand2_1 _20642_ (.A(_02390_),
    .B(_02418_),
    .Y(_02422_));
 sky130_fd_sc_hd__a21bo_1 _20643_ (.A1(_02389_),
    .A2(_02419_),
    .B1_N(_02422_),
    .X(_02423_));
 sky130_fd_sc_hd__and2_1 _20644_ (.A(_02396_),
    .B(_02401_),
    .X(_02424_));
 sky130_fd_sc_hd__a21oi_1 _20645_ (.A1(_02395_),
    .A2(_02402_),
    .B1(_02424_),
    .Y(_02425_));
 sky130_fd_sc_hd__nand2_1 _20646_ (.A(_02408_),
    .B(_02409_),
    .Y(_02426_));
 sky130_fd_sc_hd__nand2_1 _20647_ (.A(_02403_),
    .B(_02410_),
    .Y(_02427_));
 sky130_fd_sc_hd__a21bo_1 _20648_ (.A1(_02398_),
    .A2(_02400_),
    .B1_N(_02397_),
    .X(_02428_));
 sky130_fd_sc_hd__o2bb2ai_1 _20649_ (.A1_N(_02001_),
    .A2_N(_02227_),
    .B1(_02405_),
    .B2(_02406_),
    .Y(_02429_));
 sky130_fd_sc_hd__nand3_1 _20650_ (.A(_02004_),
    .B(_02016_),
    .C(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[13] ),
    .Y(_02430_));
 sky130_fd_sc_hd__a21o_1 _20651_ (.A1(_02004_),
    .A2(_02016_),
    .B1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[13] ),
    .X(_02431_));
 sky130_fd_sc_hd__nand2_1 _20652_ (.A(_02430_),
    .B(_02431_),
    .Y(_02432_));
 sky130_fd_sc_hd__nor2_1 _20653_ (.A(_02001_),
    .B(_02229_),
    .Y(_02433_));
 sky130_fd_sc_hd__xnor2_1 _20654_ (.A(_02432_),
    .B(_02433_),
    .Y(_02434_));
 sky130_fd_sc_hd__xor2_1 _20655_ (.A(_02429_),
    .B(_02434_),
    .X(_02435_));
 sky130_fd_sc_hd__xor2_1 _20656_ (.A(_02428_),
    .B(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__a21oi_1 _20657_ (.A1(_02365_),
    .A2(_02407_),
    .B1(_02364_),
    .Y(_02437_));
 sky130_fd_sc_hd__o21a_1 _20658_ (.A1(_02020_),
    .A2(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[0] ),
    .B1(_02003_),
    .X(_02438_));
 sky130_fd_sc_hd__and2b_1 _20659_ (.A_N(_02188_),
    .B(_02438_),
    .X(_02439_));
 sky130_fd_sc_hd__xnor2_2 _20660_ (.A(_02406_),
    .B(_02439_),
    .Y(_02440_));
 sky130_fd_sc_hd__xnor2_1 _20661_ (.A(_02366_),
    .B(_02440_),
    .Y(_02441_));
 sky130_fd_sc_hd__xnor2_1 _20662_ (.A(_02437_),
    .B(_02441_),
    .Y(_02442_));
 sky130_fd_sc_hd__xnor2_1 _20663_ (.A(_02436_),
    .B(_02442_),
    .Y(_02443_));
 sky130_fd_sc_hd__a21oi_1 _20664_ (.A1(_02426_),
    .A2(_02427_),
    .B1(_02443_),
    .Y(_02444_));
 sky130_fd_sc_hd__and3_1 _20665_ (.A(_02426_),
    .B(_02427_),
    .C(_02443_),
    .X(_02445_));
 sky130_fd_sc_hd__nor2_1 _20666_ (.A(_02444_),
    .B(_02445_),
    .Y(_02446_));
 sky130_fd_sc_hd__xnor2_1 _20667_ (.A(_02425_),
    .B(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__or2_1 _20668_ (.A(_02394_),
    .B(_02414_),
    .X(_02448_));
 sky130_fd_sc_hd__o21a_1 _20669_ (.A1(_02411_),
    .A2(_02413_),
    .B1(_02448_),
    .X(_02449_));
 sky130_fd_sc_hd__xor2_1 _20670_ (.A(_02447_),
    .B(_02449_),
    .X(_02450_));
 sky130_fd_sc_hd__xor2_1 _20671_ (.A(_02416_),
    .B(_02450_),
    .X(_02451_));
 sky130_fd_sc_hd__xor2_1 _20672_ (.A(_02423_),
    .B(_02451_),
    .X(_02452_));
 sky130_fd_sc_hd__or2_1 _20673_ (.A(net837),
    .B(_01386_),
    .X(_02453_));
 sky130_fd_sc_hd__o211a_1 _20674_ (.A1(_01819_),
    .A2(_02452_),
    .B1(_02453_),
    .C1(_02035_),
    .X(_00787_));
 sky130_fd_sc_hd__a21o_1 _20675_ (.A1(_02416_),
    .A2(_02422_),
    .B1(_02450_),
    .X(_02454_));
 sky130_fd_sc_hd__and2_1 _20676_ (.A(_02419_),
    .B(_02451_),
    .X(_02455_));
 sky130_fd_sc_hd__nand2_1 _20677_ (.A(_02389_),
    .B(_02455_),
    .Y(_02456_));
 sky130_fd_sc_hd__and2b_1 _20678_ (.A_N(_02449_),
    .B(_02447_),
    .X(_02457_));
 sky130_fd_sc_hd__and2_1 _20679_ (.A(_02429_),
    .B(_02434_),
    .X(_02458_));
 sky130_fd_sc_hd__a21o_1 _20680_ (.A1(_02428_),
    .A2(_02435_),
    .B1(_02458_),
    .X(_02459_));
 sky130_fd_sc_hd__nor2_1 _20681_ (.A(_02365_),
    .B(_02440_),
    .Y(_02460_));
 sky130_fd_sc_hd__and2_1 _20682_ (.A(_02364_),
    .B(_02440_),
    .X(_02461_));
 sky130_fd_sc_hd__nor2_1 _20683_ (.A(_02460_),
    .B(_02461_),
    .Y(_02462_));
 sky130_fd_sc_hd__buf_4 _20684_ (.A(_02462_),
    .X(_02463_));
 sky130_fd_sc_hd__a21bo_1 _20685_ (.A1(_02431_),
    .A2(_02433_),
    .B1_N(_02430_),
    .X(_02464_));
 sky130_fd_sc_hd__a31o_2 _20686_ (.A1(_02004_),
    .A2(_02018_),
    .A3(_02438_),
    .B1(_02227_),
    .X(_02465_));
 sky130_fd_sc_hd__buf_2 _20687_ (.A(_02465_),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_4 _20688_ (.A0(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[7] ),
    .A1(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[4] ),
    .S(_02003_),
    .X(_02467_));
 sky130_fd_sc_hd__clkbuf_4 _20689_ (.A(_02467_),
    .X(_02468_));
 sky130_fd_sc_hd__nand2_1 _20690_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[14] ),
    .B(_02468_),
    .Y(_02469_));
 sky130_fd_sc_hd__buf_2 _20691_ (.A(_02467_),
    .X(_02470_));
 sky130_fd_sc_hd__or2_1 _20692_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[14] ),
    .B(_02470_),
    .X(_02471_));
 sky130_fd_sc_hd__and3_1 _20693_ (.A(_02466_),
    .B(_02469_),
    .C(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__clkbuf_4 _20694_ (.A(_02465_),
    .X(_02473_));
 sky130_fd_sc_hd__a21oi_1 _20695_ (.A1(_02469_),
    .A2(_02471_),
    .B1(_02473_),
    .Y(_02474_));
 sky130_fd_sc_hd__nor2_1 _20696_ (.A(_02472_),
    .B(_02474_),
    .Y(_02475_));
 sky130_fd_sc_hd__xor2_1 _20697_ (.A(_02464_),
    .B(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__xnor2_1 _20698_ (.A(_02463_),
    .B(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__and2b_1 _20699_ (.A_N(_02437_),
    .B(_02441_),
    .X(_02478_));
 sky130_fd_sc_hd__a21o_1 _20700_ (.A1(_02436_),
    .A2(_02442_),
    .B1(_02478_),
    .X(_02479_));
 sky130_fd_sc_hd__and2b_1 _20701_ (.A_N(_02477_),
    .B(_02479_),
    .X(_02480_));
 sky130_fd_sc_hd__or2b_1 _20702_ (.A(_02479_),
    .B_N(_02477_),
    .X(_02481_));
 sky130_fd_sc_hd__or2b_1 _20703_ (.A(_02480_),
    .B_N(_02481_),
    .X(_02482_));
 sky130_fd_sc_hd__xnor2_1 _20704_ (.A(_02459_),
    .B(_02482_),
    .Y(_02483_));
 sky130_fd_sc_hd__o21ba_1 _20705_ (.A1(_02425_),
    .A2(_02445_),
    .B1_N(_02444_),
    .X(_02484_));
 sky130_fd_sc_hd__xnor2_1 _20706_ (.A(_02483_),
    .B(_02484_),
    .Y(_02485_));
 sky130_fd_sc_hd__xnor2_1 _20707_ (.A(_02457_),
    .B(_02485_),
    .Y(_02486_));
 sky130_fd_sc_hd__a21o_1 _20708_ (.A1(_02454_),
    .A2(_02456_),
    .B1(_02486_),
    .X(_02487_));
 sky130_fd_sc_hd__a31oi_1 _20709_ (.A1(_02486_),
    .A2(_02454_),
    .A3(_02456_),
    .B1(_06404_),
    .Y(_02488_));
 sky130_fd_sc_hd__a22o_1 _20710_ (.A1(\top_inst.deskew_buff_inst.col_input[46] ),
    .A2(_11723_),
    .B1(_02487_),
    .B2(_02488_),
    .X(_02489_));
 sky130_fd_sc_hd__and2_1 _20711_ (.A(_02135_),
    .B(_02489_),
    .X(_02490_));
 sky130_fd_sc_hd__clkbuf_1 _20712_ (.A(_02490_),
    .X(_00788_));
 sky130_fd_sc_hd__buf_4 _20713_ (.A(_06168_),
    .X(_02491_));
 sky130_fd_sc_hd__nand2_1 _20714_ (.A(_02457_),
    .B(_02485_),
    .Y(_02492_));
 sky130_fd_sc_hd__nand2_1 _20715_ (.A(_02492_),
    .B(_02487_),
    .Y(_02493_));
 sky130_fd_sc_hd__or2b_1 _20716_ (.A(_02484_),
    .B_N(_02483_),
    .X(_02494_));
 sky130_fd_sc_hd__a21oi_1 _20717_ (.A1(_02464_),
    .A2(_02475_),
    .B1(_02472_),
    .Y(_02495_));
 sky130_fd_sc_hd__nand2_1 _20718_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[15] ),
    .B(_02470_),
    .Y(_02496_));
 sky130_fd_sc_hd__or2_1 _20719_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[15] ),
    .B(_02470_),
    .X(_02497_));
 sky130_fd_sc_hd__and3_1 _20720_ (.A(_02466_),
    .B(_02496_),
    .C(_02497_),
    .X(_02498_));
 sky130_fd_sc_hd__a21oi_1 _20721_ (.A1(_02496_),
    .A2(_02497_),
    .B1(_02466_),
    .Y(_02499_));
 sky130_fd_sc_hd__nor2_1 _20722_ (.A(_02498_),
    .B(_02499_),
    .Y(_02500_));
 sky130_fd_sc_hd__xnor2_1 _20723_ (.A(_02469_),
    .B(_02500_),
    .Y(_02501_));
 sky130_fd_sc_hd__xnor2_1 _20724_ (.A(_02463_),
    .B(_02501_),
    .Y(_02502_));
 sky130_fd_sc_hd__clkbuf_4 _20725_ (.A(_02461_),
    .X(_02503_));
 sky130_fd_sc_hd__a21oi_1 _20726_ (.A1(_02463_),
    .A2(_02476_),
    .B1(_02503_),
    .Y(_02504_));
 sky130_fd_sc_hd__xnor2_1 _20727_ (.A(_02502_),
    .B(_02504_),
    .Y(_02505_));
 sky130_fd_sc_hd__xnor2_1 _20728_ (.A(_02495_),
    .B(_02505_),
    .Y(_02506_));
 sky130_fd_sc_hd__a21oi_1 _20729_ (.A1(_02459_),
    .A2(_02481_),
    .B1(_02480_),
    .Y(_02507_));
 sky130_fd_sc_hd__nor2_1 _20730_ (.A(_02506_),
    .B(_02507_),
    .Y(_02508_));
 sky130_fd_sc_hd__and2_1 _20731_ (.A(_02506_),
    .B(_02507_),
    .X(_02509_));
 sky130_fd_sc_hd__or2_1 _20732_ (.A(_02508_),
    .B(_02509_),
    .X(_02510_));
 sky130_fd_sc_hd__xnor2_2 _20733_ (.A(_02494_),
    .B(_02510_),
    .Y(_02511_));
 sky130_fd_sc_hd__nor2_1 _20734_ (.A(_02493_),
    .B(_02511_),
    .Y(_02512_));
 sky130_fd_sc_hd__a21o_1 _20735_ (.A1(_02493_),
    .A2(_02511_),
    .B1(_07595_),
    .X(_02513_));
 sky130_fd_sc_hd__o221a_1 _20736_ (.A1(net278),
    .A2(_02491_),
    .B1(_02512_),
    .B2(_02513_),
    .C1(_01863_),
    .X(_00789_));
 sky130_fd_sc_hd__nor2_1 _20737_ (.A(_02502_),
    .B(_02504_),
    .Y(_02514_));
 sky130_fd_sc_hd__nor2_1 _20738_ (.A(_02495_),
    .B(_02505_),
    .Y(_02515_));
 sky130_fd_sc_hd__o21ba_1 _20739_ (.A1(_02469_),
    .A2(_02499_),
    .B1_N(_02498_),
    .X(_02516_));
 sky130_fd_sc_hd__nand2_2 _20740_ (.A(_02364_),
    .B(_02440_),
    .Y(_02517_));
 sky130_fd_sc_hd__clkbuf_4 _20741_ (.A(_02462_),
    .X(_02518_));
 sky130_fd_sc_hd__nand2_1 _20742_ (.A(_02518_),
    .B(_02501_),
    .Y(_02519_));
 sky130_fd_sc_hd__nand2_1 _20743_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[16] ),
    .B(_02470_),
    .Y(_02520_));
 sky130_fd_sc_hd__or2_1 _20744_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[16] ),
    .B(_02467_),
    .X(_02521_));
 sky130_fd_sc_hd__and3_1 _20745_ (.A(_02465_),
    .B(_02520_),
    .C(_02521_),
    .X(_02522_));
 sky130_fd_sc_hd__a21oi_1 _20746_ (.A1(_02520_),
    .A2(_02521_),
    .B1(_02466_),
    .Y(_02523_));
 sky130_fd_sc_hd__nor2_1 _20747_ (.A(_02522_),
    .B(_02523_),
    .Y(_02524_));
 sky130_fd_sc_hd__xnor2_1 _20748_ (.A(_02496_),
    .B(_02524_),
    .Y(_02525_));
 sky130_fd_sc_hd__xnor2_1 _20749_ (.A(_02518_),
    .B(_02525_),
    .Y(_02526_));
 sky130_fd_sc_hd__a21o_1 _20750_ (.A1(_02517_),
    .A2(_02519_),
    .B1(_02526_),
    .X(_02527_));
 sky130_fd_sc_hd__clkbuf_4 _20751_ (.A(_02517_),
    .X(_02528_));
 sky130_fd_sc_hd__nand3_1 _20752_ (.A(_02528_),
    .B(_02519_),
    .C(_02526_),
    .Y(_02529_));
 sky130_fd_sc_hd__and2_1 _20753_ (.A(_02527_),
    .B(_02529_),
    .X(_02530_));
 sky130_fd_sc_hd__xnor2_1 _20754_ (.A(_02516_),
    .B(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__o21ai_2 _20755_ (.A1(_02514_),
    .A2(_02515_),
    .B1(_02531_),
    .Y(_02532_));
 sky130_fd_sc_hd__or3_1 _20756_ (.A(_02514_),
    .B(_02515_),
    .C(_02531_),
    .X(_02533_));
 sky130_fd_sc_hd__and2_1 _20757_ (.A(_02532_),
    .B(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__xnor2_1 _20758_ (.A(_02508_),
    .B(_02534_),
    .Y(_02535_));
 sky130_fd_sc_hd__nor2_1 _20759_ (.A(_02486_),
    .B(_02511_),
    .Y(_02536_));
 sky130_fd_sc_hd__nand2_1 _20760_ (.A(_02455_),
    .B(_02536_),
    .Y(_02537_));
 sky130_fd_sc_hd__a21oi_2 _20761_ (.A1(_02385_),
    .A2(_02388_),
    .B1(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__and2b_1 _20762_ (.A_N(_02454_),
    .B(_02536_),
    .X(_02539_));
 sky130_fd_sc_hd__a21oi_1 _20763_ (.A1(_02494_),
    .A2(_02492_),
    .B1(_02510_),
    .Y(_02540_));
 sky130_fd_sc_hd__nor3_1 _20764_ (.A(_02538_),
    .B(_02539_),
    .C(_02540_),
    .Y(_02541_));
 sky130_fd_sc_hd__or2_1 _20765_ (.A(_02535_),
    .B(_02541_),
    .X(_02542_));
 sky130_fd_sc_hd__nand2_1 _20766_ (.A(_02535_),
    .B(_02541_),
    .Y(_02543_));
 sky130_fd_sc_hd__and2_1 _20767_ (.A(_02542_),
    .B(_02543_),
    .X(_02544_));
 sky130_fd_sc_hd__or2_1 _20768_ (.A(net270),
    .B(_01386_),
    .X(_02545_));
 sky130_fd_sc_hd__o211a_1 _20769_ (.A1(_01819_),
    .A2(_02544_),
    .B1(_02545_),
    .C1(_02035_),
    .X(_00790_));
 sky130_fd_sc_hd__nand2_1 _20770_ (.A(_02508_),
    .B(_02534_),
    .Y(_02546_));
 sky130_fd_sc_hd__or2b_1 _20771_ (.A(_02516_),
    .B_N(_02530_),
    .X(_02547_));
 sky130_fd_sc_hd__nand2_1 _20772_ (.A(_02518_),
    .B(_02525_),
    .Y(_02548_));
 sky130_fd_sc_hd__nand2_1 _20773_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[17] ),
    .B(_02467_),
    .Y(_02549_));
 sky130_fd_sc_hd__or2_1 _20774_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[17] ),
    .B(_02467_),
    .X(_02550_));
 sky130_fd_sc_hd__and3_1 _20775_ (.A(_02465_),
    .B(_02549_),
    .C(_02550_),
    .X(_02551_));
 sky130_fd_sc_hd__a21oi_1 _20776_ (.A1(_02549_),
    .A2(_02550_),
    .B1(_02466_),
    .Y(_02552_));
 sky130_fd_sc_hd__nor2_1 _20777_ (.A(_02551_),
    .B(_02552_),
    .Y(_02553_));
 sky130_fd_sc_hd__xnor2_1 _20778_ (.A(_02520_),
    .B(_02553_),
    .Y(_02554_));
 sky130_fd_sc_hd__xnor2_1 _20779_ (.A(_02518_),
    .B(_02554_),
    .Y(_02555_));
 sky130_fd_sc_hd__a21o_1 _20780_ (.A1(_02517_),
    .A2(_02548_),
    .B1(_02555_),
    .X(_02556_));
 sky130_fd_sc_hd__nand3_1 _20781_ (.A(_02517_),
    .B(_02548_),
    .C(_02555_),
    .Y(_02557_));
 sky130_fd_sc_hd__and2_1 _20782_ (.A(_02556_),
    .B(_02557_),
    .X(_02558_));
 sky130_fd_sc_hd__clkbuf_4 _20783_ (.A(_02468_),
    .X(_02559_));
 sky130_fd_sc_hd__a31o_1 _20784_ (.A1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[15] ),
    .A2(_02559_),
    .A3(_02524_),
    .B1(_02522_),
    .X(_02560_));
 sky130_fd_sc_hd__xnor2_1 _20785_ (.A(_02558_),
    .B(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__a21o_1 _20786_ (.A1(_02527_),
    .A2(_02547_),
    .B1(_02561_),
    .X(_02562_));
 sky130_fd_sc_hd__nand3_1 _20787_ (.A(_02527_),
    .B(_02547_),
    .C(_02561_),
    .Y(_02563_));
 sky130_fd_sc_hd__nand2_1 _20788_ (.A(_02562_),
    .B(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__xor2_1 _20789_ (.A(_02532_),
    .B(_02564_),
    .X(_02565_));
 sky130_fd_sc_hd__a21oi_1 _20790_ (.A1(_02546_),
    .A2(_02542_),
    .B1(_02565_),
    .Y(_02566_));
 sky130_fd_sc_hd__a31o_1 _20791_ (.A1(_02546_),
    .A2(_02542_),
    .A3(_02565_),
    .B1(_01984_),
    .X(_02567_));
 sky130_fd_sc_hd__o221a_1 _20792_ (.A1(net280),
    .A2(_02491_),
    .B1(_02566_),
    .B2(_02567_),
    .C1(_01863_),
    .X(_00791_));
 sky130_fd_sc_hd__and2_1 _20793_ (.A(net268),
    .B(_05634_),
    .X(_02568_));
 sky130_fd_sc_hd__a21o_1 _20794_ (.A1(_02532_),
    .A2(_02546_),
    .B1(_02564_),
    .X(_02569_));
 sky130_fd_sc_hd__or2b_1 _20795_ (.A(_02535_),
    .B_N(_02565_),
    .X(_02570_));
 sky130_fd_sc_hd__or2_1 _20796_ (.A(_02541_),
    .B(_02570_),
    .X(_02571_));
 sky130_fd_sc_hd__nand2_1 _20797_ (.A(_02558_),
    .B(_02560_),
    .Y(_02572_));
 sky130_fd_sc_hd__nand2_1 _20798_ (.A(_02462_),
    .B(_02554_),
    .Y(_02573_));
 sky130_fd_sc_hd__nand2_1 _20799_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[18] ),
    .B(_02467_),
    .Y(_02574_));
 sky130_fd_sc_hd__or2_1 _20800_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[18] ),
    .B(_02467_),
    .X(_02575_));
 sky130_fd_sc_hd__and3_1 _20801_ (.A(_02465_),
    .B(_02574_),
    .C(_02575_),
    .X(_02576_));
 sky130_fd_sc_hd__a21oi_1 _20802_ (.A1(_02574_),
    .A2(_02575_),
    .B1(_02465_),
    .Y(_02577_));
 sky130_fd_sc_hd__nor2_1 _20803_ (.A(_02576_),
    .B(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__xnor2_1 _20804_ (.A(_02549_),
    .B(_02578_),
    .Y(_02579_));
 sky130_fd_sc_hd__xnor2_1 _20805_ (.A(_02462_),
    .B(_02579_),
    .Y(_02580_));
 sky130_fd_sc_hd__a21o_1 _20806_ (.A1(_02517_),
    .A2(_02573_),
    .B1(_02580_),
    .X(_02581_));
 sky130_fd_sc_hd__nand3_1 _20807_ (.A(_02517_),
    .B(_02573_),
    .C(_02580_),
    .Y(_02582_));
 sky130_fd_sc_hd__and2_1 _20808_ (.A(_02581_),
    .B(_02582_),
    .X(_02583_));
 sky130_fd_sc_hd__a31o_1 _20809_ (.A1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[16] ),
    .A2(_02559_),
    .A3(_02553_),
    .B1(_02551_),
    .X(_02584_));
 sky130_fd_sc_hd__xnor2_1 _20810_ (.A(_02583_),
    .B(_02584_),
    .Y(_02585_));
 sky130_fd_sc_hd__a21oi_2 _20811_ (.A1(_02556_),
    .A2(_02572_),
    .B1(_02585_),
    .Y(_02586_));
 sky130_fd_sc_hd__and3_1 _20812_ (.A(_02556_),
    .B(_02572_),
    .C(_02585_),
    .X(_02587_));
 sky130_fd_sc_hd__or2_1 _20813_ (.A(_02586_),
    .B(_02587_),
    .X(_02588_));
 sky130_fd_sc_hd__xnor2_1 _20814_ (.A(_02562_),
    .B(_02588_),
    .Y(_02589_));
 sky130_fd_sc_hd__a21oi_1 _20815_ (.A1(_02569_),
    .A2(_02571_),
    .B1(_02589_),
    .Y(_02590_));
 sky130_fd_sc_hd__a31o_1 _20816_ (.A1(_02589_),
    .A2(_02569_),
    .A3(_02571_),
    .B1(_05406_),
    .X(_02591_));
 sky130_fd_sc_hd__nor2_1 _20817_ (.A(_02590_),
    .B(_02591_),
    .Y(_02592_));
 sky130_fd_sc_hd__o21a_1 _20818_ (.A1(_02568_),
    .A2(_02592_),
    .B1(_04870_),
    .X(_00792_));
 sky130_fd_sc_hd__nor2_1 _20819_ (.A(_02562_),
    .B(_02588_),
    .Y(_02593_));
 sky130_fd_sc_hd__or2_1 _20820_ (.A(_02593_),
    .B(_02590_),
    .X(_02594_));
 sky130_fd_sc_hd__nand2_1 _20821_ (.A(_02463_),
    .B(_02579_),
    .Y(_02595_));
 sky130_fd_sc_hd__nand2_1 _20822_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[19] ),
    .B(_02470_),
    .Y(_02596_));
 sky130_fd_sc_hd__or2_1 _20823_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[19] ),
    .B(_02470_),
    .X(_02597_));
 sky130_fd_sc_hd__and3_1 _20824_ (.A(_02466_),
    .B(_02596_),
    .C(_02597_),
    .X(_02598_));
 sky130_fd_sc_hd__a21oi_1 _20825_ (.A1(_02596_),
    .A2(_02597_),
    .B1(_02473_),
    .Y(_02599_));
 sky130_fd_sc_hd__nor2_1 _20826_ (.A(_02598_),
    .B(_02599_),
    .Y(_02600_));
 sky130_fd_sc_hd__xnor2_1 _20827_ (.A(_02574_),
    .B(_02600_),
    .Y(_02601_));
 sky130_fd_sc_hd__xnor2_1 _20828_ (.A(_02518_),
    .B(_02601_),
    .Y(_02602_));
 sky130_fd_sc_hd__a21o_1 _20829_ (.A1(_02517_),
    .A2(_02595_),
    .B1(_02602_),
    .X(_02603_));
 sky130_fd_sc_hd__nand3_1 _20830_ (.A(_02528_),
    .B(_02595_),
    .C(_02602_),
    .Y(_02604_));
 sky130_fd_sc_hd__and2_1 _20831_ (.A(_02603_),
    .B(_02604_),
    .X(_02605_));
 sky130_fd_sc_hd__a31o_1 _20832_ (.A1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[17] ),
    .A2(_02559_),
    .A3(_02578_),
    .B1(_02576_),
    .X(_02606_));
 sky130_fd_sc_hd__xnor2_1 _20833_ (.A(_02605_),
    .B(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__nand2_1 _20834_ (.A(_02583_),
    .B(_02584_),
    .Y(_02608_));
 sky130_fd_sc_hd__nand2_1 _20835_ (.A(_02581_),
    .B(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__xor2_1 _20836_ (.A(_02607_),
    .B(_02609_),
    .X(_02610_));
 sky130_fd_sc_hd__xor2_1 _20837_ (.A(_02586_),
    .B(_02610_),
    .X(_02611_));
 sky130_fd_sc_hd__nor2_1 _20838_ (.A(_02594_),
    .B(_02611_),
    .Y(_02612_));
 sky130_fd_sc_hd__a21o_1 _20839_ (.A1(_02594_),
    .A2(_02611_),
    .B1(_07595_),
    .X(_02613_));
 sky130_fd_sc_hd__o221a_1 _20840_ (.A1(net966),
    .A2(_02491_),
    .B1(_02612_),
    .B2(_02613_),
    .C1(_01863_),
    .X(_00793_));
 sky130_fd_sc_hd__a21o_1 _20841_ (.A1(_02581_),
    .A2(_02608_),
    .B1(_02607_),
    .X(_02614_));
 sky130_fd_sc_hd__nand2_1 _20842_ (.A(_02605_),
    .B(_02606_),
    .Y(_02615_));
 sky130_fd_sc_hd__nand2_1 _20843_ (.A(_02463_),
    .B(_02601_),
    .Y(_02616_));
 sky130_fd_sc_hd__nand2_1 _20844_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[20] ),
    .B(_02468_),
    .Y(_02617_));
 sky130_fd_sc_hd__or2_1 _20845_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[20] ),
    .B(_02470_),
    .X(_02618_));
 sky130_fd_sc_hd__and3_1 _20846_ (.A(_02466_),
    .B(_02617_),
    .C(_02618_),
    .X(_02619_));
 sky130_fd_sc_hd__a21oi_1 _20847_ (.A1(_02617_),
    .A2(_02618_),
    .B1(_02473_),
    .Y(_02620_));
 sky130_fd_sc_hd__nor2_1 _20848_ (.A(_02619_),
    .B(_02620_),
    .Y(_02621_));
 sky130_fd_sc_hd__xnor2_1 _20849_ (.A(_02596_),
    .B(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__xnor2_1 _20850_ (.A(_02518_),
    .B(_02622_),
    .Y(_02623_));
 sky130_fd_sc_hd__a21o_1 _20851_ (.A1(_02517_),
    .A2(_02616_),
    .B1(_02623_),
    .X(_02624_));
 sky130_fd_sc_hd__nand3_1 _20852_ (.A(_02528_),
    .B(_02616_),
    .C(_02623_),
    .Y(_02625_));
 sky130_fd_sc_hd__and2_1 _20853_ (.A(_02624_),
    .B(_02625_),
    .X(_02626_));
 sky130_fd_sc_hd__a31o_1 _20854_ (.A1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[18] ),
    .A2(_02559_),
    .A3(_02600_),
    .B1(_02598_),
    .X(_02627_));
 sky130_fd_sc_hd__xnor2_1 _20855_ (.A(_02626_),
    .B(_02627_),
    .Y(_02628_));
 sky130_fd_sc_hd__a21o_1 _20856_ (.A1(_02603_),
    .A2(_02615_),
    .B1(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__nand3_1 _20857_ (.A(_02603_),
    .B(_02615_),
    .C(_02628_),
    .Y(_02630_));
 sky130_fd_sc_hd__nand2_1 _20858_ (.A(_02629_),
    .B(_02630_),
    .Y(_02631_));
 sky130_fd_sc_hd__xnor2_2 _20859_ (.A(_02614_),
    .B(_02631_),
    .Y(_02632_));
 sky130_fd_sc_hd__or2_1 _20860_ (.A(_02589_),
    .B(_02611_),
    .X(_02633_));
 sky130_fd_sc_hd__nor2_1 _20861_ (.A(_02586_),
    .B(_02593_),
    .Y(_02634_));
 sky130_fd_sc_hd__o22a_1 _20862_ (.A1(_02569_),
    .A2(_02633_),
    .B1(_02634_),
    .B2(_02610_),
    .X(_02635_));
 sky130_fd_sc_hd__o31a_1 _20863_ (.A1(_02541_),
    .A2(_02570_),
    .A3(_02633_),
    .B1(_02635_),
    .X(_02636_));
 sky130_fd_sc_hd__xor2_1 _20864_ (.A(_02632_),
    .B(_02636_),
    .X(_02637_));
 sky130_fd_sc_hd__clkbuf_4 _20865_ (.A(_06701_),
    .X(_02638_));
 sky130_fd_sc_hd__or2_1 _20866_ (.A(net861),
    .B(_02638_),
    .X(_02639_));
 sky130_fd_sc_hd__o211a_1 _20867_ (.A1(_01819_),
    .A2(_02637_),
    .B1(_02639_),
    .C1(_02035_),
    .X(_00794_));
 sky130_fd_sc_hd__or2_1 _20868_ (.A(_02614_),
    .B(_02631_),
    .X(_02640_));
 sky130_fd_sc_hd__o21ai_1 _20869_ (.A1(_02632_),
    .A2(_02636_),
    .B1(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__nand2_1 _20870_ (.A(_02626_),
    .B(_02627_),
    .Y(_02642_));
 sky130_fd_sc_hd__buf_4 _20871_ (.A(_02518_),
    .X(_02643_));
 sky130_fd_sc_hd__nand2_1 _20872_ (.A(_02643_),
    .B(_02622_),
    .Y(_02644_));
 sky130_fd_sc_hd__nand2_1 _20873_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[21] ),
    .B(_02468_),
    .Y(_02645_));
 sky130_fd_sc_hd__or2_1 _20874_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[21] ),
    .B(_02470_),
    .X(_02646_));
 sky130_fd_sc_hd__nand2_1 _20875_ (.A(_02645_),
    .B(_02646_),
    .Y(_02647_));
 sky130_fd_sc_hd__xnor2_2 _20876_ (.A(_02473_),
    .B(_02647_),
    .Y(_02648_));
 sky130_fd_sc_hd__xnor2_1 _20877_ (.A(_02617_),
    .B(_02648_),
    .Y(_02649_));
 sky130_fd_sc_hd__xnor2_1 _20878_ (.A(_02463_),
    .B(_02649_),
    .Y(_02650_));
 sky130_fd_sc_hd__a21o_1 _20879_ (.A1(_02528_),
    .A2(_02644_),
    .B1(_02650_),
    .X(_02651_));
 sky130_fd_sc_hd__nand3_1 _20880_ (.A(_02528_),
    .B(_02644_),
    .C(_02650_),
    .Y(_02652_));
 sky130_fd_sc_hd__and2_1 _20881_ (.A(_02651_),
    .B(_02652_),
    .X(_02653_));
 sky130_fd_sc_hd__a31o_1 _20882_ (.A1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[19] ),
    .A2(_02559_),
    .A3(_02621_),
    .B1(_02619_),
    .X(_02654_));
 sky130_fd_sc_hd__xnor2_1 _20883_ (.A(_02653_),
    .B(_02654_),
    .Y(_02655_));
 sky130_fd_sc_hd__a21o_1 _20884_ (.A1(_02624_),
    .A2(_02642_),
    .B1(_02655_),
    .X(_02656_));
 sky130_fd_sc_hd__nand3_1 _20885_ (.A(_02624_),
    .B(_02642_),
    .C(_02655_),
    .Y(_02657_));
 sky130_fd_sc_hd__nand2_1 _20886_ (.A(_02656_),
    .B(_02657_),
    .Y(_02658_));
 sky130_fd_sc_hd__xnor2_1 _20887_ (.A(_02629_),
    .B(_02658_),
    .Y(_02659_));
 sky130_fd_sc_hd__xnor2_1 _20888_ (.A(_02641_),
    .B(_02659_),
    .Y(_02660_));
 sky130_fd_sc_hd__or2_1 _20889_ (.A(net782),
    .B(_02638_),
    .X(_02661_));
 sky130_fd_sc_hd__o211a_1 _20890_ (.A1(_01819_),
    .A2(_02660_),
    .B1(_02661_),
    .C1(_02035_),
    .X(_00795_));
 sky130_fd_sc_hd__or2_1 _20891_ (.A(_02632_),
    .B(_02659_),
    .X(_02662_));
 sky130_fd_sc_hd__a21o_1 _20892_ (.A1(_02629_),
    .A2(_02640_),
    .B1(_02658_),
    .X(_02663_));
 sky130_fd_sc_hd__o21a_1 _20893_ (.A1(_02636_),
    .A2(_02662_),
    .B1(_02663_),
    .X(_02664_));
 sky130_fd_sc_hd__nand2_1 _20894_ (.A(_02653_),
    .B(_02654_),
    .Y(_02665_));
 sky130_fd_sc_hd__or2_1 _20895_ (.A(_02466_),
    .B(_02468_),
    .X(_02666_));
 sky130_fd_sc_hd__nand2_1 _20896_ (.A(_02473_),
    .B(_02646_),
    .Y(_02667_));
 sky130_fd_sc_hd__o21a_1 _20897_ (.A1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[21] ),
    .A2(_02666_),
    .B1(_02667_),
    .X(_02668_));
 sky130_fd_sc_hd__xnor2_1 _20898_ (.A(_02518_),
    .B(_02668_),
    .Y(_02669_));
 sky130_fd_sc_hd__a21o_1 _20899_ (.A1(_02463_),
    .A2(_02649_),
    .B1(_02503_),
    .X(_02670_));
 sky130_fd_sc_hd__or2b_1 _20900_ (.A(_02669_),
    .B_N(_02670_),
    .X(_02671_));
 sky130_fd_sc_hd__or2b_1 _20901_ (.A(_02670_),
    .B_N(_02669_),
    .X(_02672_));
 sky130_fd_sc_hd__nand2_1 _20902_ (.A(_02671_),
    .B(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hd__a31oi_4 _20903_ (.A1(_02004_),
    .A2(_02018_),
    .A3(_02438_),
    .B1(_02227_),
    .Y(_02674_));
 sky130_fd_sc_hd__nor2_1 _20904_ (.A(_02674_),
    .B(_02647_),
    .Y(_02675_));
 sky130_fd_sc_hd__a31oi_2 _20905_ (.A1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[20] ),
    .A2(_02559_),
    .A3(_02648_),
    .B1(_02675_),
    .Y(_02676_));
 sky130_fd_sc_hd__xnor2_1 _20906_ (.A(_02673_),
    .B(_02676_),
    .Y(_02677_));
 sky130_fd_sc_hd__a21oi_2 _20907_ (.A1(_02651_),
    .A2(_02665_),
    .B1(_02677_),
    .Y(_02678_));
 sky130_fd_sc_hd__and3_1 _20908_ (.A(_02651_),
    .B(_02665_),
    .C(_02677_),
    .X(_02679_));
 sky130_fd_sc_hd__or2_1 _20909_ (.A(_02678_),
    .B(_02679_),
    .X(_02680_));
 sky130_fd_sc_hd__xnor2_1 _20910_ (.A(_02656_),
    .B(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__nor2_1 _20911_ (.A(_05405_),
    .B(_02681_),
    .Y(_02682_));
 sky130_fd_sc_hd__a22o_1 _20912_ (.A1(\top_inst.deskew_buff_inst.col_input[54] ),
    .A2(_11723_),
    .B1(_02664_),
    .B2(_02682_),
    .X(_02683_));
 sky130_fd_sc_hd__and2_1 _20913_ (.A(_02135_),
    .B(_02683_),
    .X(_02684_));
 sky130_fd_sc_hd__clkbuf_1 _20914_ (.A(_02684_),
    .X(_00796_));
 sky130_fd_sc_hd__nor2_1 _20915_ (.A(_02656_),
    .B(_02680_),
    .Y(_02685_));
 sky130_fd_sc_hd__or2b_1 _20916_ (.A(_02685_),
    .B_N(_02664_),
    .X(_02686_));
 sky130_fd_sc_hd__and2_1 _20917_ (.A(_02518_),
    .B(_02668_),
    .X(_02687_));
 sky130_fd_sc_hd__nand2_1 _20918_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[23] ),
    .B(_02470_),
    .Y(_02688_));
 sky130_fd_sc_hd__or2_1 _20919_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[23] ),
    .B(_02467_),
    .X(_02689_));
 sky130_fd_sc_hd__and3_1 _20920_ (.A(_02465_),
    .B(_02688_),
    .C(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__a21oi_1 _20921_ (.A1(_02688_),
    .A2(_02689_),
    .B1(_02466_),
    .Y(_02691_));
 sky130_fd_sc_hd__nor2_1 _20922_ (.A(_02690_),
    .B(_02691_),
    .Y(_02692_));
 sky130_fd_sc_hd__xnor2_1 _20923_ (.A(_02645_),
    .B(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__xor2_1 _20924_ (.A(_02518_),
    .B(_02693_),
    .X(_02694_));
 sky130_fd_sc_hd__o21ai_1 _20925_ (.A1(_02503_),
    .A2(_02687_),
    .B1(_02694_),
    .Y(_02695_));
 sky130_fd_sc_hd__or3_1 _20926_ (.A(_02503_),
    .B(_02687_),
    .C(_02694_),
    .X(_02696_));
 sky130_fd_sc_hd__nand2_1 _20927_ (.A(_02695_),
    .B(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__or2_1 _20928_ (.A(_02667_),
    .B(_02697_),
    .X(_02698_));
 sky130_fd_sc_hd__nand2_1 _20929_ (.A(_02667_),
    .B(_02697_),
    .Y(_02699_));
 sky130_fd_sc_hd__and2_1 _20930_ (.A(_02698_),
    .B(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__o21a_1 _20931_ (.A1(_02673_),
    .A2(_02676_),
    .B1(_02671_),
    .X(_02701_));
 sky130_fd_sc_hd__xnor2_1 _20932_ (.A(_02700_),
    .B(_02701_),
    .Y(_02702_));
 sky130_fd_sc_hd__xor2_1 _20933_ (.A(_02678_),
    .B(_02702_),
    .X(_02703_));
 sky130_fd_sc_hd__xor2_1 _20934_ (.A(_02686_),
    .B(_02703_),
    .X(_02704_));
 sky130_fd_sc_hd__or2_1 _20935_ (.A(net647),
    .B(_02638_),
    .X(_02705_));
 sky130_fd_sc_hd__buf_6 _20936_ (.A(_04868_),
    .X(_02706_));
 sky130_fd_sc_hd__buf_4 _20937_ (.A(_02706_),
    .X(_02707_));
 sky130_fd_sc_hd__o211a_1 _20938_ (.A1(_01819_),
    .A2(_02704_),
    .B1(_02705_),
    .C1(_02707_),
    .X(_00797_));
 sky130_fd_sc_hd__or2b_1 _20939_ (.A(_02681_),
    .B_N(_02703_),
    .X(_02708_));
 sky130_fd_sc_hd__nor2_1 _20940_ (.A(_02662_),
    .B(_02708_),
    .Y(_02709_));
 sky130_fd_sc_hd__and2b_1 _20941_ (.A_N(_02635_),
    .B(_02709_),
    .X(_02710_));
 sky130_fd_sc_hd__nor2_1 _20942_ (.A(_02570_),
    .B(_02633_),
    .Y(_02711_));
 sky130_fd_sc_hd__o311a_1 _20943_ (.A1(_02538_),
    .A2(_02539_),
    .A3(_02540_),
    .B1(_02711_),
    .C1(_02709_),
    .X(_02712_));
 sky130_fd_sc_hd__o21ai_1 _20944_ (.A1(_02678_),
    .A2(_02685_),
    .B1(_02702_),
    .Y(_02713_));
 sky130_fd_sc_hd__o21ai_1 _20945_ (.A1(_02663_),
    .A2(_02708_),
    .B1(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__nor3_1 _20946_ (.A(_02710_),
    .B(_02712_),
    .C(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__or2b_1 _20947_ (.A(_02701_),
    .B_N(_02700_),
    .X(_02716_));
 sky130_fd_sc_hd__nand2_1 _20948_ (.A(_02643_),
    .B(_02693_),
    .Y(_02717_));
 sky130_fd_sc_hd__nand2_1 _20949_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[24] ),
    .B(_02468_),
    .Y(_02718_));
 sky130_fd_sc_hd__or2_1 _20950_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[24] ),
    .B(_02468_),
    .X(_02719_));
 sky130_fd_sc_hd__and3_1 _20951_ (.A(_02473_),
    .B(_02718_),
    .C(_02719_),
    .X(_02720_));
 sky130_fd_sc_hd__a21oi_1 _20952_ (.A1(_02718_),
    .A2(_02719_),
    .B1(_02473_),
    .Y(_02721_));
 sky130_fd_sc_hd__nor2_1 _20953_ (.A(_02720_),
    .B(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__xnor2_1 _20954_ (.A(_02688_),
    .B(_02722_),
    .Y(_02723_));
 sky130_fd_sc_hd__xnor2_1 _20955_ (.A(_02643_),
    .B(_02723_),
    .Y(_02724_));
 sky130_fd_sc_hd__a21o_1 _20956_ (.A1(_02528_),
    .A2(_02717_),
    .B1(_02724_),
    .X(_02725_));
 sky130_fd_sc_hd__nand3_1 _20957_ (.A(_02528_),
    .B(_02717_),
    .C(_02724_),
    .Y(_02726_));
 sky130_fd_sc_hd__and2_1 _20958_ (.A(_02725_),
    .B(_02726_),
    .X(_02727_));
 sky130_fd_sc_hd__a31o_1 _20959_ (.A1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[21] ),
    .A2(_02559_),
    .A3(_02692_),
    .B1(_02690_),
    .X(_02728_));
 sky130_fd_sc_hd__xnor2_1 _20960_ (.A(_02727_),
    .B(_02728_),
    .Y(_02729_));
 sky130_fd_sc_hd__a21o_1 _20961_ (.A1(_02695_),
    .A2(_02698_),
    .B1(_02729_),
    .X(_02730_));
 sky130_fd_sc_hd__nand3_1 _20962_ (.A(_02695_),
    .B(_02698_),
    .C(_02729_),
    .Y(_02731_));
 sky130_fd_sc_hd__nand2_1 _20963_ (.A(_02730_),
    .B(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__or2_2 _20964_ (.A(_02716_),
    .B(_02732_),
    .X(_02733_));
 sky130_fd_sc_hd__nand2_1 _20965_ (.A(_02716_),
    .B(_02732_),
    .Y(_02734_));
 sky130_fd_sc_hd__nand2_1 _20966_ (.A(_02733_),
    .B(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__or2_1 _20967_ (.A(_02715_),
    .B(_02735_),
    .X(_02736_));
 sky130_fd_sc_hd__nand2_1 _20968_ (.A(_02715_),
    .B(_02735_),
    .Y(_02737_));
 sky130_fd_sc_hd__and2_1 _20969_ (.A(_02736_),
    .B(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__or2_1 _20970_ (.A(net696),
    .B(_02638_),
    .X(_02739_));
 sky130_fd_sc_hd__o211a_1 _20971_ (.A1(_01819_),
    .A2(_02738_),
    .B1(_02739_),
    .C1(_02707_),
    .X(_00798_));
 sky130_fd_sc_hd__nand2_1 _20972_ (.A(_02727_),
    .B(_02728_),
    .Y(_02740_));
 sky130_fd_sc_hd__nand2_1 _20973_ (.A(_02643_),
    .B(_02723_),
    .Y(_02741_));
 sky130_fd_sc_hd__nand2_1 _20974_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[25] ),
    .B(_02468_),
    .Y(_02742_));
 sky130_fd_sc_hd__or2_1 _20975_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[25] ),
    .B(_02470_),
    .X(_02743_));
 sky130_fd_sc_hd__and3_1 _20976_ (.A(_02466_),
    .B(_02742_),
    .C(_02743_),
    .X(_02744_));
 sky130_fd_sc_hd__a21oi_1 _20977_ (.A1(_02742_),
    .A2(_02743_),
    .B1(_02473_),
    .Y(_02745_));
 sky130_fd_sc_hd__nor2_1 _20978_ (.A(_02744_),
    .B(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__xnor2_1 _20979_ (.A(_02718_),
    .B(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__xnor2_1 _20980_ (.A(_02463_),
    .B(_02747_),
    .Y(_02748_));
 sky130_fd_sc_hd__a21o_1 _20981_ (.A1(_02528_),
    .A2(_02741_),
    .B1(_02748_),
    .X(_02749_));
 sky130_fd_sc_hd__nand3_1 _20982_ (.A(_02528_),
    .B(_02741_),
    .C(_02748_),
    .Y(_02750_));
 sky130_fd_sc_hd__and2_1 _20983_ (.A(_02749_),
    .B(_02750_),
    .X(_02751_));
 sky130_fd_sc_hd__a31o_1 _20984_ (.A1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[23] ),
    .A2(_02559_),
    .A3(_02722_),
    .B1(_02720_),
    .X(_02752_));
 sky130_fd_sc_hd__xnor2_1 _20985_ (.A(_02751_),
    .B(_02752_),
    .Y(_02753_));
 sky130_fd_sc_hd__a21o_1 _20986_ (.A1(_02725_),
    .A2(_02740_),
    .B1(_02753_),
    .X(_02754_));
 sky130_fd_sc_hd__nand3_1 _20987_ (.A(_02725_),
    .B(_02740_),
    .C(_02753_),
    .Y(_02755_));
 sky130_fd_sc_hd__nand2_1 _20988_ (.A(_02754_),
    .B(_02755_),
    .Y(_02756_));
 sky130_fd_sc_hd__xor2_1 _20989_ (.A(_02730_),
    .B(_02756_),
    .X(_02757_));
 sky130_fd_sc_hd__a21oi_1 _20990_ (.A1(_02733_),
    .A2(_02736_),
    .B1(_02757_),
    .Y(_02758_));
 sky130_fd_sc_hd__a31o_1 _20991_ (.A1(_02733_),
    .A2(_02736_),
    .A3(_02757_),
    .B1(_01984_),
    .X(_02759_));
 sky130_fd_sc_hd__o221a_1 _20992_ (.A1(net919),
    .A2(_02491_),
    .B1(_02758_),
    .B2(_02759_),
    .C1(_01863_),
    .X(_00799_));
 sky130_fd_sc_hd__or2b_1 _20993_ (.A(_02735_),
    .B_N(_02757_),
    .X(_02760_));
 sky130_fd_sc_hd__a21oi_1 _20994_ (.A1(_02730_),
    .A2(_02733_),
    .B1(_02756_),
    .Y(_02761_));
 sky130_fd_sc_hd__inv_2 _20995_ (.A(_02761_),
    .Y(_02762_));
 sky130_fd_sc_hd__o21a_1 _20996_ (.A1(_02715_),
    .A2(_02760_),
    .B1(_02762_),
    .X(_02763_));
 sky130_fd_sc_hd__nand2_1 _20997_ (.A(_02751_),
    .B(_02752_),
    .Y(_02764_));
 sky130_fd_sc_hd__nand2_1 _20998_ (.A(_02473_),
    .B(_02743_),
    .Y(_02765_));
 sky130_fd_sc_hd__o21a_1 _20999_ (.A1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[25] ),
    .A2(_02666_),
    .B1(_02765_),
    .X(_02766_));
 sky130_fd_sc_hd__xnor2_1 _21000_ (.A(_02463_),
    .B(_02766_),
    .Y(_02767_));
 sky130_fd_sc_hd__a21o_1 _21001_ (.A1(_02463_),
    .A2(_02747_),
    .B1(_02503_),
    .X(_02768_));
 sky130_fd_sc_hd__or2b_1 _21002_ (.A(_02767_),
    .B_N(_02768_),
    .X(_02769_));
 sky130_fd_sc_hd__or2b_1 _21003_ (.A(_02768_),
    .B_N(_02767_),
    .X(_02770_));
 sky130_fd_sc_hd__nand2_1 _21004_ (.A(_02769_),
    .B(_02770_),
    .Y(_02771_));
 sky130_fd_sc_hd__o21ba_1 _21005_ (.A1(_02718_),
    .A2(_02745_),
    .B1_N(_02744_),
    .X(_02772_));
 sky130_fd_sc_hd__xnor2_1 _21006_ (.A(_02771_),
    .B(_02772_),
    .Y(_02773_));
 sky130_fd_sc_hd__a21oi_2 _21007_ (.A1(_02749_),
    .A2(_02764_),
    .B1(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__and3_1 _21008_ (.A(_02749_),
    .B(_02764_),
    .C(_02773_),
    .X(_02775_));
 sky130_fd_sc_hd__or2_1 _21009_ (.A(_02774_),
    .B(_02775_),
    .X(_02776_));
 sky130_fd_sc_hd__and2_1 _21010_ (.A(_02754_),
    .B(_02776_),
    .X(_02777_));
 sky130_fd_sc_hd__nor2_1 _21011_ (.A(_02754_),
    .B(_02776_),
    .Y(_02778_));
 sky130_fd_sc_hd__or2_1 _21012_ (.A(_02777_),
    .B(_02778_),
    .X(_02779_));
 sky130_fd_sc_hd__nor2_1 _21013_ (.A(_05405_),
    .B(_02779_),
    .Y(_02780_));
 sky130_fd_sc_hd__a22o_1 _21014_ (.A1(\top_inst.deskew_buff_inst.col_input[58] ),
    .A2(_11723_),
    .B1(_02763_),
    .B2(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__and2_1 _21015_ (.A(_02135_),
    .B(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__clkbuf_1 _21016_ (.A(_02782_),
    .X(_00800_));
 sky130_fd_sc_hd__inv_2 _21017_ (.A(_02778_),
    .Y(_02783_));
 sky130_fd_sc_hd__inv_2 _21018_ (.A(_02765_),
    .Y(_02784_));
 sky130_fd_sc_hd__and2_1 _21019_ (.A(_02643_),
    .B(_02766_),
    .X(_02785_));
 sky130_fd_sc_hd__nand2_2 _21020_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[27] ),
    .B(_02468_),
    .Y(_02786_));
 sky130_fd_sc_hd__or2_1 _21021_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[27] ),
    .B(_02468_),
    .X(_02787_));
 sky130_fd_sc_hd__nand2_1 _21022_ (.A(_02786_),
    .B(_02787_),
    .Y(_02788_));
 sky130_fd_sc_hd__xnor2_1 _21023_ (.A(_02473_),
    .B(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__a21oi_1 _21024_ (.A1(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[25] ),
    .A2(_02559_),
    .B1(_02789_),
    .Y(_02790_));
 sky130_fd_sc_hd__and3_1 _21025_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[25] ),
    .B(_02559_),
    .C(_02789_),
    .X(_02791_));
 sky130_fd_sc_hd__nor2_1 _21026_ (.A(_02790_),
    .B(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__xor2_2 _21027_ (.A(_02643_),
    .B(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__o21ai_2 _21028_ (.A1(_02503_),
    .A2(_02785_),
    .B1(_02793_),
    .Y(_02794_));
 sky130_fd_sc_hd__or3_1 _21029_ (.A(_02503_),
    .B(_02785_),
    .C(_02793_),
    .X(_02795_));
 sky130_fd_sc_hd__nand3_1 _21030_ (.A(_02784_),
    .B(_02794_),
    .C(_02795_),
    .Y(_02796_));
 sky130_fd_sc_hd__a21o_1 _21031_ (.A1(_02794_),
    .A2(_02795_),
    .B1(_02784_),
    .X(_02797_));
 sky130_fd_sc_hd__and2_1 _21032_ (.A(_02796_),
    .B(_02797_),
    .X(_02798_));
 sky130_fd_sc_hd__o21a_1 _21033_ (.A1(_02771_),
    .A2(_02772_),
    .B1(_02769_),
    .X(_02799_));
 sky130_fd_sc_hd__xnor2_2 _21034_ (.A(_02798_),
    .B(_02799_),
    .Y(_02800_));
 sky130_fd_sc_hd__xor2_1 _21035_ (.A(_02774_),
    .B(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__and3_1 _21036_ (.A(_02763_),
    .B(_02783_),
    .C(_02801_),
    .X(_02802_));
 sky130_fd_sc_hd__a21o_1 _21037_ (.A1(_02763_),
    .A2(_02783_),
    .B1(_02801_),
    .X(_02803_));
 sky130_fd_sc_hd__nand2_1 _21038_ (.A(_06178_),
    .B(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__o221a_1 _21039_ (.A1(net997),
    .A2(_02491_),
    .B1(_02802_),
    .B2(_02804_),
    .C1(_01863_),
    .X(_00801_));
 sky130_fd_sc_hd__or2b_1 _21040_ (.A(_02779_),
    .B_N(_02801_),
    .X(_02805_));
 sky130_fd_sc_hd__nor2_1 _21041_ (.A(_02760_),
    .B(_02805_),
    .Y(_02806_));
 sky130_fd_sc_hd__o31ai_2 _21042_ (.A1(_02710_),
    .A2(_02712_),
    .A3(_02714_),
    .B1(_02806_),
    .Y(_02807_));
 sky130_fd_sc_hd__o21ai_1 _21043_ (.A1(_02774_),
    .A2(_02778_),
    .B1(_02800_),
    .Y(_02808_));
 sky130_fd_sc_hd__o21a_1 _21044_ (.A1(_02762_),
    .A2(_02805_),
    .B1(_02808_),
    .X(_02809_));
 sky130_fd_sc_hd__or2b_1 _21045_ (.A(_02799_),
    .B_N(_02798_),
    .X(_02810_));
 sky130_fd_sc_hd__xnor2_1 _21046_ (.A(_02746_),
    .B(_02786_),
    .Y(_02811_));
 sky130_fd_sc_hd__and2_1 _21047_ (.A(_02643_),
    .B(_02811_),
    .X(_02812_));
 sky130_fd_sc_hd__nor2_1 _21048_ (.A(_02643_),
    .B(_02811_),
    .Y(_02813_));
 sky130_fd_sc_hd__or2_1 _21049_ (.A(_02812_),
    .B(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__a21oi_2 _21050_ (.A1(_02643_),
    .A2(_02792_),
    .B1(_02503_),
    .Y(_02815_));
 sky130_fd_sc_hd__or2_1 _21051_ (.A(_02814_),
    .B(_02815_),
    .X(_02816_));
 sky130_fd_sc_hd__nand2_1 _21052_ (.A(_02814_),
    .B(_02815_),
    .Y(_02817_));
 sky130_fd_sc_hd__nand2_1 _21053_ (.A(_02816_),
    .B(_02817_),
    .Y(_02818_));
 sky130_fd_sc_hd__o21ba_1 _21054_ (.A1(_02674_),
    .A2(_02788_),
    .B1_N(_02791_),
    .X(_02819_));
 sky130_fd_sc_hd__xnor2_1 _21055_ (.A(_02818_),
    .B(_02819_),
    .Y(_02820_));
 sky130_fd_sc_hd__a21oi_1 _21056_ (.A1(_02794_),
    .A2(_02796_),
    .B1(_02820_),
    .Y(_02821_));
 sky130_fd_sc_hd__and3_1 _21057_ (.A(_02794_),
    .B(_02796_),
    .C(_02820_),
    .X(_02822_));
 sky130_fd_sc_hd__or2_1 _21058_ (.A(_02821_),
    .B(_02822_),
    .X(_02823_));
 sky130_fd_sc_hd__and2_1 _21059_ (.A(_02810_),
    .B(_02823_),
    .X(_02824_));
 sky130_fd_sc_hd__nor2_1 _21060_ (.A(_02810_),
    .B(_02823_),
    .Y(_02825_));
 sky130_fd_sc_hd__or2_1 _21061_ (.A(_02824_),
    .B(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__a21oi_2 _21062_ (.A1(_02807_),
    .A2(_02809_),
    .B1(_02826_),
    .Y(_02827_));
 sky130_fd_sc_hd__and3_1 _21063_ (.A(_02807_),
    .B(_02809_),
    .C(_02826_),
    .X(_02828_));
 sky130_fd_sc_hd__o21ai_1 _21064_ (.A1(_02827_),
    .A2(_02828_),
    .B1(_06178_),
    .Y(_02829_));
 sky130_fd_sc_hd__o211a_1 _21065_ (.A1(net869),
    .A2(_01735_),
    .B1(_02829_),
    .C1(_02707_),
    .X(_00802_));
 sky130_fd_sc_hd__o21ai_1 _21066_ (.A1(_02503_),
    .A2(_02812_),
    .B1(_02793_),
    .Y(_02830_));
 sky130_fd_sc_hd__or3_1 _21067_ (.A(_02503_),
    .B(_02793_),
    .C(_02812_),
    .X(_02831_));
 sky130_fd_sc_hd__nand2_1 _21068_ (.A(_02830_),
    .B(_02831_),
    .Y(_02832_));
 sky130_fd_sc_hd__o21ba_1 _21069_ (.A1(_02745_),
    .A2(_02786_),
    .B1_N(_02744_),
    .X(_02833_));
 sky130_fd_sc_hd__xor2_1 _21070_ (.A(_02832_),
    .B(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__o21a_1 _21071_ (.A1(_02818_),
    .A2(_02819_),
    .B1(_02816_),
    .X(_02835_));
 sky130_fd_sc_hd__xnor2_1 _21072_ (.A(_02834_),
    .B(_02835_),
    .Y(_02836_));
 sky130_fd_sc_hd__xnor2_1 _21073_ (.A(_02821_),
    .B(_02836_),
    .Y(_02837_));
 sky130_fd_sc_hd__o21a_1 _21074_ (.A1(_02825_),
    .A2(net228),
    .B1(_02837_),
    .X(_02838_));
 sky130_fd_sc_hd__o31ai_2 _21075_ (.A1(_02825_),
    .A2(_02827_),
    .A3(_02837_),
    .B1(_05313_),
    .Y(_02839_));
 sky130_fd_sc_hd__o221a_1 _21076_ (.A1(net327),
    .A2(_02491_),
    .B1(_02838_),
    .B2(_02839_),
    .C1(_01863_),
    .X(_00803_));
 sky130_fd_sc_hd__or2b_1 _21077_ (.A(_02835_),
    .B_N(_02834_),
    .X(_02840_));
 sky130_fd_sc_hd__mux2_1 _21078_ (.A0(_02674_),
    .A1(_02789_),
    .S(_02786_),
    .X(_02841_));
 sky130_fd_sc_hd__xnor2_1 _21079_ (.A(_02643_),
    .B(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__xor2_1 _21080_ (.A(_02815_),
    .B(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__xnor2_1 _21081_ (.A(_02819_),
    .B(_02843_),
    .Y(_02844_));
 sky130_fd_sc_hd__inv_2 _21082_ (.A(_02844_),
    .Y(_02845_));
 sky130_fd_sc_hd__o21a_1 _21083_ (.A1(_02832_),
    .A2(_02833_),
    .B1(_02830_),
    .X(_02846_));
 sky130_fd_sc_hd__xnor2_1 _21084_ (.A(_02845_),
    .B(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__o21a_1 _21085_ (.A1(_02821_),
    .A2(_02825_),
    .B1(_02836_),
    .X(_02848_));
 sky130_fd_sc_hd__nor2_1 _21086_ (.A(_02827_),
    .B(_02848_),
    .Y(_02849_));
 sky130_fd_sc_hd__o21a_1 _21087_ (.A1(_02840_),
    .A2(_02847_),
    .B1(_02849_),
    .X(_02850_));
 sky130_fd_sc_hd__a21oi_1 _21088_ (.A1(_02840_),
    .A2(_02847_),
    .B1(_05406_),
    .Y(_02851_));
 sky130_fd_sc_hd__a22oi_1 _21089_ (.A1(net1097),
    .A2(_05328_),
    .B1(_02850_),
    .B2(_02851_),
    .Y(_02852_));
 sky130_fd_sc_hd__nor2_1 _21090_ (.A(_05440_),
    .B(_02852_),
    .Y(_00804_));
 sky130_fd_sc_hd__or2b_1 _21091_ (.A(_02819_),
    .B_N(_02843_),
    .X(_02853_));
 sky130_fd_sc_hd__o221a_1 _21092_ (.A1(_02815_),
    .A2(_02842_),
    .B1(_02845_),
    .B2(_02846_),
    .C1(_02853_),
    .X(_02854_));
 sky130_fd_sc_hd__o21a_1 _21093_ (.A1(_02460_),
    .A2(_02841_),
    .B1(_02528_),
    .X(_02855_));
 sky130_fd_sc_hd__xnor2_1 _21094_ (.A(_02854_),
    .B(_02855_),
    .Y(_02856_));
 sky130_fd_sc_hd__xnor2_1 _21095_ (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[31] ),
    .B(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__and2b_1 _21096_ (.A_N(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[27] ),
    .B(_02666_),
    .X(_02858_));
 sky130_fd_sc_hd__xnor2_1 _21097_ (.A(_02857_),
    .B(_02858_),
    .Y(_02859_));
 sky130_fd_sc_hd__xnor2_1 _21098_ (.A(_02850_),
    .B(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__nor2_1 _21099_ (.A(net1102),
    .B(_05313_),
    .Y(_02861_));
 sky130_fd_sc_hd__a211oi_1 _21100_ (.A1(_05317_),
    .A2(_02860_),
    .B1(_02861_),
    .C1(_04867_),
    .Y(_00805_));
 sky130_fd_sc_hd__clkbuf_4 _21101_ (.A(\top_inst.grid_inst.data_path_wires[17][0] ),
    .X(_02862_));
 sky130_fd_sc_hd__or2_1 _21102_ (.A(_02862_),
    .B(_11133_),
    .X(_02863_));
 sky130_fd_sc_hd__o211a_1 _21103_ (.A1(_01987_),
    .A2(_11142_),
    .B1(_02863_),
    .C1(_02707_),
    .X(_00806_));
 sky130_fd_sc_hd__clkbuf_4 _21104_ (.A(\top_inst.grid_inst.data_path_wires[17][1] ),
    .X(_02864_));
 sky130_fd_sc_hd__or2_1 _21105_ (.A(_02864_),
    .B(_11133_),
    .X(_02865_));
 sky130_fd_sc_hd__o211a_1 _21106_ (.A1(_01990_),
    .A2(_11142_),
    .B1(_02865_),
    .C1(_02707_),
    .X(_00807_));
 sky130_fd_sc_hd__clkbuf_4 _21107_ (.A(\top_inst.grid_inst.data_path_wires[17][2] ),
    .X(_02866_));
 sky130_fd_sc_hd__or2_1 _21108_ (.A(_02866_),
    .B(_11133_),
    .X(_02867_));
 sky130_fd_sc_hd__o211a_1 _21109_ (.A1(_01993_),
    .A2(_11142_),
    .B1(_02867_),
    .C1(_02707_),
    .X(_00808_));
 sky130_fd_sc_hd__clkbuf_4 _21110_ (.A(\top_inst.grid_inst.data_path_wires[17][3] ),
    .X(_02868_));
 sky130_fd_sc_hd__buf_2 _21111_ (.A(_06619_),
    .X(_02869_));
 sky130_fd_sc_hd__or2_1 _21112_ (.A(_02868_),
    .B(_02869_),
    .X(_02870_));
 sky130_fd_sc_hd__o211a_1 _21113_ (.A1(_01995_),
    .A2(_11142_),
    .B1(_02870_),
    .C1(_02707_),
    .X(_00809_));
 sky130_fd_sc_hd__clkbuf_4 _21114_ (.A(\top_inst.grid_inst.data_path_wires[17][4] ),
    .X(_02871_));
 sky130_fd_sc_hd__or2_1 _21115_ (.A(_02871_),
    .B(_02869_),
    .X(_02872_));
 sky130_fd_sc_hd__o211a_1 _21116_ (.A1(_01997_),
    .A2(_11142_),
    .B1(_02872_),
    .C1(_02707_),
    .X(_00810_));
 sky130_fd_sc_hd__clkbuf_4 _21117_ (.A(\top_inst.grid_inst.data_path_wires[17][5] ),
    .X(_02873_));
 sky130_fd_sc_hd__or2_1 _21118_ (.A(_02873_),
    .B(_02869_),
    .X(_02874_));
 sky130_fd_sc_hd__o211a_1 _21119_ (.A1(_01999_),
    .A2(_11142_),
    .B1(_02874_),
    .C1(_02707_),
    .X(_00811_));
 sky130_fd_sc_hd__clkbuf_4 _21120_ (.A(\top_inst.grid_inst.data_path_wires[17][6] ),
    .X(_02875_));
 sky130_fd_sc_hd__or2_1 _21121_ (.A(_02875_),
    .B(_02869_),
    .X(_02876_));
 sky130_fd_sc_hd__o211a_1 _21122_ (.A1(_02001_),
    .A2(_11142_),
    .B1(_02876_),
    .C1(_02707_),
    .X(_00812_));
 sky130_fd_sc_hd__clkbuf_8 _21123_ (.A(_10583_),
    .X(_02877_));
 sky130_fd_sc_hd__clkbuf_4 _21124_ (.A(\top_inst.grid_inst.data_path_wires[17][7] ),
    .X(_02878_));
 sky130_fd_sc_hd__or2_1 _21125_ (.A(_02878_),
    .B(_02869_),
    .X(_02879_));
 sky130_fd_sc_hd__clkbuf_4 _21126_ (.A(_02706_),
    .X(_02880_));
 sky130_fd_sc_hd__o211a_1 _21127_ (.A1(_02004_),
    .A2(_02877_),
    .B1(_02879_),
    .C1(_02880_),
    .X(_00813_));
 sky130_fd_sc_hd__clkbuf_4 _21128_ (.A(_05269_),
    .X(_02881_));
 sky130_fd_sc_hd__clkbuf_4 _21129_ (.A(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[0] ),
    .X(_02882_));
 sky130_fd_sc_hd__clkbuf_4 _21130_ (.A(_02882_),
    .X(_02883_));
 sky130_fd_sc_hd__or2_1 _21131_ (.A(_02883_),
    .B(_02021_),
    .X(_02884_));
 sky130_fd_sc_hd__o211a_1 _21132_ (.A1(_02862_),
    .A2(_02881_),
    .B1(_02884_),
    .C1(_02880_),
    .X(_00814_));
 sky130_fd_sc_hd__clkbuf_4 _21133_ (.A(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[1] ),
    .X(_02885_));
 sky130_fd_sc_hd__or2_1 _21134_ (.A(_02885_),
    .B(_02021_),
    .X(_02886_));
 sky130_fd_sc_hd__o211a_1 _21135_ (.A1(_02864_),
    .A2(_02881_),
    .B1(_02886_),
    .C1(_02880_),
    .X(_00815_));
 sky130_fd_sc_hd__clkbuf_4 _21136_ (.A(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[2] ),
    .X(_02887_));
 sky130_fd_sc_hd__or2_1 _21137_ (.A(_02887_),
    .B(_02021_),
    .X(_02888_));
 sky130_fd_sc_hd__o211a_1 _21138_ (.A1(_02866_),
    .A2(_02881_),
    .B1(_02888_),
    .C1(_02880_),
    .X(_00816_));
 sky130_fd_sc_hd__buf_2 _21139_ (.A(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[3] ),
    .X(_02889_));
 sky130_fd_sc_hd__or2_1 _21140_ (.A(_02889_),
    .B(_02021_),
    .X(_02890_));
 sky130_fd_sc_hd__o211a_1 _21141_ (.A1(_02868_),
    .A2(_02881_),
    .B1(_02890_),
    .C1(_02880_),
    .X(_00817_));
 sky130_fd_sc_hd__clkbuf_4 _21142_ (.A(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[4] ),
    .X(_02891_));
 sky130_fd_sc_hd__or2_1 _21143_ (.A(_02891_),
    .B(_02021_),
    .X(_02892_));
 sky130_fd_sc_hd__o211a_1 _21144_ (.A1(_02871_),
    .A2(_02881_),
    .B1(_02892_),
    .C1(_02880_),
    .X(_00818_));
 sky130_fd_sc_hd__buf_2 _21145_ (.A(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[5] ),
    .X(_02893_));
 sky130_fd_sc_hd__or2_1 _21146_ (.A(_02893_),
    .B(_02021_),
    .X(_02894_));
 sky130_fd_sc_hd__o211a_1 _21147_ (.A1(_02873_),
    .A2(_02881_),
    .B1(_02894_),
    .C1(_02880_),
    .X(_00819_));
 sky130_fd_sc_hd__buf_2 _21148_ (.A(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[6] ),
    .X(_02895_));
 sky130_fd_sc_hd__or2_1 _21149_ (.A(_02895_),
    .B(_02021_),
    .X(_02896_));
 sky130_fd_sc_hd__o211a_1 _21150_ (.A1(_02875_),
    .A2(_02881_),
    .B1(_02896_),
    .C1(_02880_),
    .X(_00820_));
 sky130_fd_sc_hd__clkbuf_4 _21151_ (.A(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[7] ),
    .X(_02897_));
 sky130_fd_sc_hd__or2_1 _21152_ (.A(_02897_),
    .B(_02021_),
    .X(_02898_));
 sky130_fd_sc_hd__o211a_1 _21153_ (.A1(_02878_),
    .A2(_02881_),
    .B1(_02898_),
    .C1(_02880_),
    .X(_00821_));
 sky130_fd_sc_hd__and3_1 _21154_ (.A(_02862_),
    .B(_02883_),
    .C(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[0] ),
    .X(_02899_));
 sky130_fd_sc_hd__a21oi_1 _21155_ (.A1(_02862_),
    .A2(_02883_),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[0] ),
    .Y(_02900_));
 sky130_fd_sc_hd__o21ai_1 _21156_ (.A1(_02899_),
    .A2(_02900_),
    .B1(_06178_),
    .Y(_02901_));
 sky130_fd_sc_hd__o211a_1 _21157_ (.A1(net454),
    .A2(_01735_),
    .B1(_02901_),
    .C1(_02880_),
    .X(_00822_));
 sky130_fd_sc_hd__a22o_1 _21158_ (.A1(\top_inst.grid_inst.data_path_wires[17][0] ),
    .A2(_02885_),
    .B1(_02883_),
    .B2(_02864_),
    .X(_02902_));
 sky130_fd_sc_hd__nand4_2 _21159_ (.A(_02864_),
    .B(_02862_),
    .C(_02885_),
    .D(_02883_),
    .Y(_02903_));
 sky130_fd_sc_hd__nand3_1 _21160_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[1] ),
    .B(_02902_),
    .C(_02903_),
    .Y(_02904_));
 sky130_fd_sc_hd__a21o_1 _21161_ (.A1(_02902_),
    .A2(_02903_),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[1] ),
    .X(_02905_));
 sky130_fd_sc_hd__a21o_1 _21162_ (.A1(_02904_),
    .A2(_02905_),
    .B1(_02899_),
    .X(_02906_));
 sky130_fd_sc_hd__nand3_2 _21163_ (.A(_02899_),
    .B(_02904_),
    .C(_02905_),
    .Y(_02907_));
 sky130_fd_sc_hd__a21o_1 _21164_ (.A1(_02906_),
    .A2(_02907_),
    .B1(_05732_),
    .X(_02908_));
 sky130_fd_sc_hd__clkbuf_4 _21165_ (.A(_02706_),
    .X(_02909_));
 sky130_fd_sc_hd__o211a_1 _21166_ (.A1(net325),
    .A2(_06169_),
    .B1(_02908_),
    .C1(_02909_),
    .X(_00823_));
 sky130_fd_sc_hd__nand2_1 _21167_ (.A(_02862_),
    .B(_02887_),
    .Y(_02910_));
 sky130_fd_sc_hd__a22o_1 _21168_ (.A1(_02864_),
    .A2(_02885_),
    .B1(_02883_),
    .B2(_02866_),
    .X(_02911_));
 sky130_fd_sc_hd__nand4_1 _21169_ (.A(_02866_),
    .B(_02864_),
    .C(_02885_),
    .D(_02883_),
    .Y(_02912_));
 sky130_fd_sc_hd__nand2_1 _21170_ (.A(_02911_),
    .B(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__xor2_1 _21171_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[2] ),
    .B(_02913_),
    .X(_02914_));
 sky130_fd_sc_hd__nand2_1 _21172_ (.A(_02903_),
    .B(_02904_),
    .Y(_02915_));
 sky130_fd_sc_hd__xor2_1 _21173_ (.A(_02914_),
    .B(_02915_),
    .X(_02916_));
 sky130_fd_sc_hd__or2_1 _21174_ (.A(_02910_),
    .B(_02916_),
    .X(_02917_));
 sky130_fd_sc_hd__nand2_1 _21175_ (.A(_02910_),
    .B(_02916_),
    .Y(_02918_));
 sky130_fd_sc_hd__and2_1 _21176_ (.A(_02917_),
    .B(_02918_),
    .X(_02919_));
 sky130_fd_sc_hd__xnor2_1 _21177_ (.A(_02907_),
    .B(_02919_),
    .Y(_02920_));
 sky130_fd_sc_hd__or2_1 _21178_ (.A(net282),
    .B(_02638_),
    .X(_02921_));
 sky130_fd_sc_hd__o211a_1 _21179_ (.A1(_01819_),
    .A2(_02920_),
    .B1(_02921_),
    .C1(_02909_),
    .X(_00824_));
 sky130_fd_sc_hd__or2b_1 _21180_ (.A(_02907_),
    .B_N(_02919_),
    .X(_02922_));
 sky130_fd_sc_hd__or2b_1 _21181_ (.A(_02914_),
    .B_N(_02915_),
    .X(_02923_));
 sky130_fd_sc_hd__a22o_1 _21182_ (.A1(_02862_),
    .A2(_02889_),
    .B1(_02887_),
    .B2(_02864_),
    .X(_02924_));
 sky130_fd_sc_hd__and3_1 _21183_ (.A(\top_inst.grid_inst.data_path_wires[17][1] ),
    .B(\top_inst.grid_inst.data_path_wires[17][0] ),
    .C(_02889_),
    .X(_02925_));
 sky130_fd_sc_hd__nand2_2 _21184_ (.A(_02887_),
    .B(_02925_),
    .Y(_02926_));
 sky130_fd_sc_hd__nand2_1 _21185_ (.A(_02924_),
    .B(_02926_),
    .Y(_02927_));
 sky130_fd_sc_hd__a22o_1 _21186_ (.A1(_02866_),
    .A2(_02885_),
    .B1(_02882_),
    .B2(_02868_),
    .X(_02928_));
 sky130_fd_sc_hd__nand4_1 _21187_ (.A(_02868_),
    .B(_02866_),
    .C(_02885_),
    .D(_02883_),
    .Y(_02929_));
 sky130_fd_sc_hd__and3_1 _21188_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[3] ),
    .B(_02928_),
    .C(_02929_),
    .X(_02930_));
 sky130_fd_sc_hd__a21oi_1 _21189_ (.A1(_02928_),
    .A2(_02929_),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[3] ),
    .Y(_02931_));
 sky130_fd_sc_hd__or2_1 _21190_ (.A(_02930_),
    .B(_02931_),
    .X(_02932_));
 sky130_fd_sc_hd__a21boi_2 _21191_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[2] ),
    .A2(_02911_),
    .B1_N(_02912_),
    .Y(_02933_));
 sky130_fd_sc_hd__xnor2_1 _21192_ (.A(_02932_),
    .B(_02933_),
    .Y(_02934_));
 sky130_fd_sc_hd__xnor2_1 _21193_ (.A(_02927_),
    .B(_02934_),
    .Y(_02935_));
 sky130_fd_sc_hd__a21o_1 _21194_ (.A1(_02923_),
    .A2(_02917_),
    .B1(_02935_),
    .X(_02936_));
 sky130_fd_sc_hd__inv_2 _21195_ (.A(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__and3_1 _21196_ (.A(_02923_),
    .B(_02917_),
    .C(_02935_),
    .X(_02938_));
 sky130_fd_sc_hd__or3_1 _21197_ (.A(_02922_),
    .B(_02937_),
    .C(_02938_),
    .X(_02939_));
 sky130_fd_sc_hd__o21ai_1 _21198_ (.A1(_02937_),
    .A2(_02938_),
    .B1(_02922_),
    .Y(_02940_));
 sky130_fd_sc_hd__and2_1 _21199_ (.A(\top_inst.deskew_buff_inst.col_input[67] ),
    .B(_05730_),
    .X(_02941_));
 sky130_fd_sc_hd__a31o_1 _21200_ (.A1(_05312_),
    .A2(_02939_),
    .A3(_02940_),
    .B1(_02941_),
    .X(_02942_));
 sky130_fd_sc_hd__and2_1 _21201_ (.A(_02135_),
    .B(_02942_),
    .X(_02943_));
 sky130_fd_sc_hd__clkbuf_1 _21202_ (.A(_02943_),
    .X(_00825_));
 sky130_fd_sc_hd__a22o_1 _21203_ (.A1(\top_inst.grid_inst.data_path_wires[17][3] ),
    .A2(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[1] ),
    .B1(_02882_),
    .B2(\top_inst.grid_inst.data_path_wires[17][4] ),
    .X(_02944_));
 sky130_fd_sc_hd__nand4_1 _21204_ (.A(_02871_),
    .B(_02868_),
    .C(_02885_),
    .D(_02882_),
    .Y(_02945_));
 sky130_fd_sc_hd__nand2_1 _21205_ (.A(_02944_),
    .B(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__xor2_2 _21206_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[4] ),
    .B(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__xor2_2 _21207_ (.A(_02926_),
    .B(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__a21bo_1 _21208_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[3] ),
    .A2(_02928_),
    .B1_N(_02929_),
    .X(_02949_));
 sky130_fd_sc_hd__xnor2_2 _21209_ (.A(_02948_),
    .B(_02949_),
    .Y(_02950_));
 sky130_fd_sc_hd__nand2_1 _21210_ (.A(_02866_),
    .B(_02887_),
    .Y(_02951_));
 sky130_fd_sc_hd__a22o_1 _21211_ (.A1(\top_inst.grid_inst.data_path_wires[17][0] ),
    .A2(_02891_),
    .B1(_02889_),
    .B2(\top_inst.grid_inst.data_path_wires[17][1] ),
    .X(_02952_));
 sky130_fd_sc_hd__a21bo_1 _21212_ (.A1(_02891_),
    .A2(_02925_),
    .B1_N(_02952_),
    .X(_02953_));
 sky130_fd_sc_hd__xor2_2 _21213_ (.A(_02951_),
    .B(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__xor2_2 _21214_ (.A(_02950_),
    .B(_02954_),
    .X(_02955_));
 sky130_fd_sc_hd__or2_1 _21215_ (.A(_02927_),
    .B(_02934_),
    .X(_02956_));
 sky130_fd_sc_hd__o21ai_2 _21216_ (.A1(_02932_),
    .A2(_02933_),
    .B1(_02956_),
    .Y(_02957_));
 sky130_fd_sc_hd__xor2_2 _21217_ (.A(_02955_),
    .B(_02957_),
    .X(_02958_));
 sky130_fd_sc_hd__nand2_1 _21218_ (.A(_02936_),
    .B(_02939_),
    .Y(_02959_));
 sky130_fd_sc_hd__nor2_1 _21219_ (.A(_02958_),
    .B(_02959_),
    .Y(_02960_));
 sky130_fd_sc_hd__a21o_1 _21220_ (.A1(_02958_),
    .A2(_02959_),
    .B1(_07595_),
    .X(_02961_));
 sky130_fd_sc_hd__buf_4 _21221_ (.A(_07707_),
    .X(_02962_));
 sky130_fd_sc_hd__o221a_1 _21222_ (.A1(net604),
    .A2(_02491_),
    .B1(_02960_),
    .B2(_02961_),
    .C1(_02962_),
    .X(_00826_));
 sky130_fd_sc_hd__nor2_1 _21223_ (.A(_02939_),
    .B(_02958_),
    .Y(_02963_));
 sky130_fd_sc_hd__and2b_1 _21224_ (.A_N(_02950_),
    .B(_02954_),
    .X(_02964_));
 sky130_fd_sc_hd__nand2_1 _21225_ (.A(_02862_),
    .B(_02893_),
    .Y(_02965_));
 sky130_fd_sc_hd__nand2_1 _21226_ (.A(_02868_),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[2] ),
    .Y(_02966_));
 sky130_fd_sc_hd__and3_1 _21227_ (.A(\top_inst.grid_inst.data_path_wires[17][2] ),
    .B(\top_inst.grid_inst.data_path_wires[17][1] ),
    .C(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[4] ),
    .X(_02967_));
 sky130_fd_sc_hd__a22o_1 _21228_ (.A1(\top_inst.grid_inst.data_path_wires[17][1] ),
    .A2(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[17][2] ),
    .X(_02968_));
 sky130_fd_sc_hd__a21bo_1 _21229_ (.A1(_02889_),
    .A2(_02967_),
    .B1_N(_02968_),
    .X(_02969_));
 sky130_fd_sc_hd__xor2_2 _21230_ (.A(_02966_),
    .B(_02969_),
    .X(_02970_));
 sky130_fd_sc_hd__xnor2_2 _21231_ (.A(_02965_),
    .B(_02970_),
    .Y(_02971_));
 sky130_fd_sc_hd__a21boi_2 _21232_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[4] ),
    .A2(_02944_),
    .B1_N(_02945_),
    .Y(_02972_));
 sky130_fd_sc_hd__a32o_1 _21233_ (.A1(_02866_),
    .A2(_02887_),
    .A3(_02952_),
    .B1(_02925_),
    .B2(_02891_),
    .X(_02973_));
 sky130_fd_sc_hd__a22o_1 _21234_ (.A1(\top_inst.grid_inst.data_path_wires[17][4] ),
    .A2(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[1] ),
    .B1(_02882_),
    .B2(\top_inst.grid_inst.data_path_wires[17][5] ),
    .X(_02974_));
 sky130_fd_sc_hd__nand4_1 _21235_ (.A(_02873_),
    .B(\top_inst.grid_inst.data_path_wires[17][4] ),
    .C(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[1] ),
    .D(_02882_),
    .Y(_02975_));
 sky130_fd_sc_hd__nand2_1 _21236_ (.A(_02974_),
    .B(_02975_),
    .Y(_02976_));
 sky130_fd_sc_hd__xor2_2 _21237_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[5] ),
    .B(_02976_),
    .X(_02977_));
 sky130_fd_sc_hd__xnor2_2 _21238_ (.A(_02973_),
    .B(_02977_),
    .Y(_02978_));
 sky130_fd_sc_hd__xnor2_2 _21239_ (.A(_02972_),
    .B(_02978_),
    .Y(_02979_));
 sky130_fd_sc_hd__xor2_2 _21240_ (.A(_02971_),
    .B(_02979_),
    .X(_02980_));
 sky130_fd_sc_hd__xor2_2 _21241_ (.A(_02964_),
    .B(_02980_),
    .X(_02981_));
 sky130_fd_sc_hd__nor2_1 _21242_ (.A(_02926_),
    .B(_02947_),
    .Y(_02982_));
 sky130_fd_sc_hd__a21o_1 _21243_ (.A1(_02948_),
    .A2(_02949_),
    .B1(_02982_),
    .X(_02983_));
 sky130_fd_sc_hd__xnor2_2 _21244_ (.A(_02981_),
    .B(_02983_),
    .Y(_02984_));
 sky130_fd_sc_hd__or2b_1 _21245_ (.A(_02955_),
    .B_N(_02957_),
    .X(_02985_));
 sky130_fd_sc_hd__o21a_1 _21246_ (.A1(_02936_),
    .A2(_02958_),
    .B1(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__xor2_1 _21247_ (.A(_02984_),
    .B(_02986_),
    .X(_02987_));
 sky130_fd_sc_hd__nand2_1 _21248_ (.A(_02963_),
    .B(_02987_),
    .Y(_02988_));
 sky130_fd_sc_hd__o21a_1 _21249_ (.A1(_02963_),
    .A2(_02987_),
    .B1(_10831_),
    .X(_02989_));
 sky130_fd_sc_hd__a22o_1 _21250_ (.A1(\top_inst.deskew_buff_inst.col_input[69] ),
    .A2(_11723_),
    .B1(_02988_),
    .B2(_02989_),
    .X(_02990_));
 sky130_fd_sc_hd__and2_1 _21251_ (.A(_02135_),
    .B(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__clkbuf_1 _21252_ (.A(_02991_),
    .X(_00827_));
 sky130_fd_sc_hd__nor2_1 _21253_ (.A(_02985_),
    .B(_02984_),
    .Y(_02992_));
 sky130_fd_sc_hd__nand2_1 _21254_ (.A(_02964_),
    .B(_02980_),
    .Y(_02993_));
 sky130_fd_sc_hd__nand2_1 _21255_ (.A(_02981_),
    .B(_02983_),
    .Y(_02994_));
 sky130_fd_sc_hd__or2b_1 _21256_ (.A(_02977_),
    .B_N(_02973_),
    .X(_02995_));
 sky130_fd_sc_hd__or2b_1 _21257_ (.A(_02972_),
    .B_N(_02978_),
    .X(_02996_));
 sky130_fd_sc_hd__and2_1 _21258_ (.A(_02971_),
    .B(_02979_),
    .X(_02997_));
 sky130_fd_sc_hd__a21boi_1 _21259_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[5] ),
    .A2(_02974_),
    .B1_N(_02975_),
    .Y(_02998_));
 sky130_fd_sc_hd__o2bb2a_1 _21260_ (.A1_N(_02889_),
    .A2_N(_02967_),
    .B1(_02969_),
    .B2(_02966_),
    .X(_02999_));
 sky130_fd_sc_hd__a22o_1 _21261_ (.A1(\top_inst.grid_inst.data_path_wires[17][5] ),
    .A2(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[1] ),
    .B1(_02882_),
    .B2(\top_inst.grid_inst.data_path_wires[17][6] ),
    .X(_03000_));
 sky130_fd_sc_hd__nand4_1 _21262_ (.A(\top_inst.grid_inst.data_path_wires[17][6] ),
    .B(\top_inst.grid_inst.data_path_wires[17][5] ),
    .C(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[1] ),
    .D(_02882_),
    .Y(_03001_));
 sky130_fd_sc_hd__and3_1 _21263_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[6] ),
    .B(_03000_),
    .C(_03001_),
    .X(_03002_));
 sky130_fd_sc_hd__a21oi_1 _21264_ (.A1(_03000_),
    .A2(_03001_),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[6] ),
    .Y(_03003_));
 sky130_fd_sc_hd__or2_1 _21265_ (.A(_03002_),
    .B(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__xor2_1 _21266_ (.A(_02999_),
    .B(_03004_),
    .X(_03005_));
 sky130_fd_sc_hd__xnor2_1 _21267_ (.A(_02998_),
    .B(_03005_),
    .Y(_03006_));
 sky130_fd_sc_hd__or2b_1 _21268_ (.A(_02965_),
    .B_N(_02970_),
    .X(_03007_));
 sky130_fd_sc_hd__a22oi_1 _21269_ (.A1(_02862_),
    .A2(_02895_),
    .B1(_02893_),
    .B2(_02864_),
    .Y(_03008_));
 sky130_fd_sc_hd__and4_1 _21270_ (.A(_02864_),
    .B(\top_inst.grid_inst.data_path_wires[17][0] ),
    .C(_02895_),
    .D(_02893_),
    .X(_03009_));
 sky130_fd_sc_hd__nor2_1 _21271_ (.A(_03008_),
    .B(_03009_),
    .Y(_03010_));
 sky130_fd_sc_hd__a22oi_1 _21272_ (.A1(\top_inst.grid_inst.data_path_wires[17][2] ),
    .A2(_02891_),
    .B1(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[17][3] ),
    .Y(_03011_));
 sky130_fd_sc_hd__and4_1 _21273_ (.A(\top_inst.grid_inst.data_path_wires[17][3] ),
    .B(\top_inst.grid_inst.data_path_wires[17][2] ),
    .C(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[3] ),
    .X(_03012_));
 sky130_fd_sc_hd__and4bb_1 _21274_ (.A_N(_03011_),
    .B_N(_03012_),
    .C(_02871_),
    .D(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[2] ),
    .X(_03013_));
 sky130_fd_sc_hd__o2bb2a_1 _21275_ (.A1_N(_02871_),
    .A2_N(_02887_),
    .B1(_03011_),
    .B2(_03012_),
    .X(_03014_));
 sky130_fd_sc_hd__nor2_1 _21276_ (.A(_03013_),
    .B(_03014_),
    .Y(_03015_));
 sky130_fd_sc_hd__xnor2_1 _21277_ (.A(_03010_),
    .B(_03015_),
    .Y(_03016_));
 sky130_fd_sc_hd__xor2_1 _21278_ (.A(_03007_),
    .B(_03016_),
    .X(_03017_));
 sky130_fd_sc_hd__nand2_1 _21279_ (.A(_03006_),
    .B(_03017_),
    .Y(_03018_));
 sky130_fd_sc_hd__or2_1 _21280_ (.A(_03006_),
    .B(_03017_),
    .X(_03019_));
 sky130_fd_sc_hd__and3_1 _21281_ (.A(_02997_),
    .B(_03018_),
    .C(_03019_),
    .X(_03020_));
 sky130_fd_sc_hd__a21oi_1 _21282_ (.A1(_03018_),
    .A2(_03019_),
    .B1(_02997_),
    .Y(_03021_));
 sky130_fd_sc_hd__a211oi_2 _21283_ (.A1(_02995_),
    .A2(_02996_),
    .B1(_03020_),
    .C1(_03021_),
    .Y(_03022_));
 sky130_fd_sc_hd__o211a_1 _21284_ (.A1(_03020_),
    .A2(_03021_),
    .B1(_02995_),
    .C1(_02996_),
    .X(_03023_));
 sky130_fd_sc_hd__a211o_1 _21285_ (.A1(_02993_),
    .A2(_02994_),
    .B1(_03022_),
    .C1(_03023_),
    .X(_03024_));
 sky130_fd_sc_hd__o211ai_1 _21286_ (.A1(_03022_),
    .A2(_03023_),
    .B1(_02993_),
    .C1(_02994_),
    .Y(_03025_));
 sky130_fd_sc_hd__and3_1 _21287_ (.A(_02992_),
    .B(_03024_),
    .C(_03025_),
    .X(_03026_));
 sky130_fd_sc_hd__a21oi_1 _21288_ (.A1(_03024_),
    .A2(_03025_),
    .B1(_02992_),
    .Y(_03027_));
 sky130_fd_sc_hd__nor2_1 _21289_ (.A(_03026_),
    .B(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__o31a_1 _21290_ (.A1(_02936_),
    .A2(_02958_),
    .A3(_02984_),
    .B1(_02988_),
    .X(_03029_));
 sky130_fd_sc_hd__xnor2_1 _21291_ (.A(_03028_),
    .B(_03029_),
    .Y(_03030_));
 sky130_fd_sc_hd__mux2_1 _21292_ (.A0(\top_inst.deskew_buff_inst.col_input[70] ),
    .A1(_03030_),
    .S(_06140_),
    .X(_03031_));
 sky130_fd_sc_hd__and2_1 _21293_ (.A(_02135_),
    .B(_03031_),
    .X(_03032_));
 sky130_fd_sc_hd__clkbuf_1 _21294_ (.A(_03032_),
    .X(_00828_));
 sky130_fd_sc_hd__or2b_1 _21295_ (.A(_02998_),
    .B_N(_03005_),
    .X(_03033_));
 sky130_fd_sc_hd__o21ai_1 _21296_ (.A1(_02999_),
    .A2(_03004_),
    .B1(_03033_),
    .Y(_03034_));
 sky130_fd_sc_hd__o21ai_1 _21297_ (.A1(_03007_),
    .A2(_03016_),
    .B1(_03018_),
    .Y(_03035_));
 sky130_fd_sc_hd__a21bo_1 _21298_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[6] ),
    .A2(_03000_),
    .B1_N(_03001_),
    .X(_03036_));
 sky130_fd_sc_hd__nor2_1 _21299_ (.A(_03012_),
    .B(_03013_),
    .Y(_03037_));
 sky130_fd_sc_hd__a22o_1 _21300_ (.A1(_02875_),
    .A2(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[1] ),
    .B1(_02882_),
    .B2(_02878_),
    .X(_03038_));
 sky130_fd_sc_hd__nand4_1 _21301_ (.A(_02878_),
    .B(_02875_),
    .C(_02885_),
    .D(_02883_),
    .Y(_03039_));
 sky130_fd_sc_hd__nand2_1 _21302_ (.A(_03038_),
    .B(_03039_),
    .Y(_03040_));
 sky130_fd_sc_hd__xor2_2 _21303_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[7] ),
    .B(_03040_),
    .X(_03041_));
 sky130_fd_sc_hd__xor2_2 _21304_ (.A(_03037_),
    .B(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__xnor2_2 _21305_ (.A(_03036_),
    .B(_03042_),
    .Y(_03043_));
 sky130_fd_sc_hd__and2_1 _21306_ (.A(_03010_),
    .B(_03015_),
    .X(_03044_));
 sky130_fd_sc_hd__a22o_1 _21307_ (.A1(\top_inst.grid_inst.data_path_wires[17][3] ),
    .A2(_02891_),
    .B1(_02889_),
    .B2(\top_inst.grid_inst.data_path_wires[17][4] ),
    .X(_03045_));
 sky130_fd_sc_hd__nand4_1 _21308_ (.A(_02871_),
    .B(_02868_),
    .C(_02891_),
    .D(_02889_),
    .Y(_03046_));
 sky130_fd_sc_hd__nand2_1 _21309_ (.A(_03045_),
    .B(_03046_),
    .Y(_03047_));
 sky130_fd_sc_hd__and2_1 _21310_ (.A(_02873_),
    .B(_02887_),
    .X(_03048_));
 sky130_fd_sc_hd__xor2_1 _21311_ (.A(_03047_),
    .B(_03048_),
    .X(_03049_));
 sky130_fd_sc_hd__nand2_1 _21312_ (.A(\top_inst.grid_inst.data_path_wires[17][2] ),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[5] ),
    .Y(_03050_));
 sky130_fd_sc_hd__nand2_1 _21313_ (.A(\top_inst.grid_inst.data_path_wires[17][1] ),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[6] ),
    .Y(_03051_));
 sky130_fd_sc_hd__and2b_1 _21314_ (.A_N(\top_inst.grid_inst.data_path_wires[17][0] ),
    .B(_02897_),
    .X(_03052_));
 sky130_fd_sc_hd__xnor2_1 _21315_ (.A(_03051_),
    .B(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__xnor2_1 _21316_ (.A(_03050_),
    .B(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__xnor2_1 _21317_ (.A(_03009_),
    .B(_03054_),
    .Y(_03055_));
 sky130_fd_sc_hd__xor2_1 _21318_ (.A(_03049_),
    .B(_03055_),
    .X(_03056_));
 sky130_fd_sc_hd__xnor2_1 _21319_ (.A(_03044_),
    .B(_03056_),
    .Y(_03057_));
 sky130_fd_sc_hd__xnor2_1 _21320_ (.A(_03043_),
    .B(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__xor2_1 _21321_ (.A(_03035_),
    .B(_03058_),
    .X(_03059_));
 sky130_fd_sc_hd__xnor2_1 _21322_ (.A(_03034_),
    .B(_03059_),
    .Y(_03060_));
 sky130_fd_sc_hd__nor2_1 _21323_ (.A(_03020_),
    .B(_03022_),
    .Y(_03061_));
 sky130_fd_sc_hd__xnor2_1 _21324_ (.A(_03060_),
    .B(_03061_),
    .Y(_03062_));
 sky130_fd_sc_hd__xnor2_1 _21325_ (.A(_02897_),
    .B(_03062_),
    .Y(_03063_));
 sky130_fd_sc_hd__xor2_1 _21326_ (.A(_03024_),
    .B(_03063_),
    .X(_03064_));
 sky130_fd_sc_hd__o21bai_1 _21327_ (.A1(_03027_),
    .A2(_03029_),
    .B1_N(_03026_),
    .Y(_03065_));
 sky130_fd_sc_hd__nor2_1 _21328_ (.A(_03064_),
    .B(_03065_),
    .Y(_03066_));
 sky130_fd_sc_hd__a21o_1 _21329_ (.A1(_03064_),
    .A2(_03065_),
    .B1(_05353_),
    .X(_03067_));
 sky130_fd_sc_hd__a2bb2o_1 _21330_ (.A1_N(_03066_),
    .A2_N(_03067_),
    .B1(\top_inst.deskew_buff_inst.col_input[71] ),
    .B2(_05354_),
    .X(_03068_));
 sky130_fd_sc_hd__and2_1 _21331_ (.A(_02135_),
    .B(_03068_),
    .X(_03069_));
 sky130_fd_sc_hd__clkbuf_1 _21332_ (.A(_03069_),
    .X(_00829_));
 sky130_fd_sc_hd__buf_4 _21333_ (.A(_07057_),
    .X(_03070_));
 sky130_fd_sc_hd__nor2_1 _21334_ (.A(_03024_),
    .B(_03063_),
    .Y(_03071_));
 sky130_fd_sc_hd__a21o_2 _21335_ (.A1(_03064_),
    .A2(_03065_),
    .B1(_03071_),
    .X(_03072_));
 sky130_fd_sc_hd__nor2_1 _21336_ (.A(_03037_),
    .B(_03041_),
    .Y(_03073_));
 sky130_fd_sc_hd__a21o_1 _21337_ (.A1(_03036_),
    .A2(_03042_),
    .B1(_03073_),
    .X(_03074_));
 sky130_fd_sc_hd__a21boi_2 _21338_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[7] ),
    .A2(_03038_),
    .B1_N(_03039_),
    .Y(_03075_));
 sky130_fd_sc_hd__a21boi_2 _21339_ (.A1(_03045_),
    .A2(_03048_),
    .B1_N(_03046_),
    .Y(_03076_));
 sky130_fd_sc_hd__and3_1 _21340_ (.A(\top_inst.grid_inst.data_path_wires[17][7] ),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[1] ),
    .C(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[0] ),
    .X(_03077_));
 sky130_fd_sc_hd__o21ai_2 _21341_ (.A1(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[1] ),
    .A2(_02882_),
    .B1(\top_inst.grid_inst.data_path_wires[17][7] ),
    .Y(_03078_));
 sky130_fd_sc_hd__nor2_1 _21342_ (.A(_03077_),
    .B(_03078_),
    .Y(_03079_));
 sky130_fd_sc_hd__buf_4 _21343_ (.A(_03079_),
    .X(_03080_));
 sky130_fd_sc_hd__xnor2_2 _21344_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[8] ),
    .B(_03080_),
    .Y(_03081_));
 sky130_fd_sc_hd__xor2_2 _21345_ (.A(_03076_),
    .B(_03081_),
    .X(_03082_));
 sky130_fd_sc_hd__xnor2_2 _21346_ (.A(_03075_),
    .B(_03082_),
    .Y(_03083_));
 sky130_fd_sc_hd__a22o_1 _21347_ (.A1(_02871_),
    .A2(_02891_),
    .B1(_02889_),
    .B2(_02873_),
    .X(_03084_));
 sky130_fd_sc_hd__nand4_1 _21348_ (.A(_02873_),
    .B(_02871_),
    .C(_02891_),
    .D(_02889_),
    .Y(_03085_));
 sky130_fd_sc_hd__nand2_1 _21349_ (.A(_03084_),
    .B(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__and2_1 _21350_ (.A(_02875_),
    .B(_02887_),
    .X(_03087_));
 sky130_fd_sc_hd__xnor2_2 _21351_ (.A(_03086_),
    .B(_03087_),
    .Y(_03088_));
 sky130_fd_sc_hd__nand2_1 _21352_ (.A(_02868_),
    .B(_02893_),
    .Y(_03089_));
 sky130_fd_sc_hd__and2b_1 _21353_ (.A_N(\top_inst.grid_inst.data_path_wires[17][1] ),
    .B(_02897_),
    .X(_03090_));
 sky130_fd_sc_hd__nand2_1 _21354_ (.A(\top_inst.grid_inst.data_path_wires[17][2] ),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[6] ),
    .Y(_03091_));
 sky130_fd_sc_hd__xnor2_2 _21355_ (.A(_03090_),
    .B(_03091_),
    .Y(_03092_));
 sky130_fd_sc_hd__xnor2_2 _21356_ (.A(_03089_),
    .B(_03092_),
    .Y(_03093_));
 sky130_fd_sc_hd__and3_1 _21357_ (.A(\top_inst.grid_inst.data_path_wires[17][1] ),
    .B(_02895_),
    .C(_03052_),
    .X(_03094_));
 sky130_fd_sc_hd__a31o_1 _21358_ (.A1(_02866_),
    .A2(_02893_),
    .A3(_03053_),
    .B1(_03094_),
    .X(_03095_));
 sky130_fd_sc_hd__xor2_2 _21359_ (.A(_03093_),
    .B(_03095_),
    .X(_03096_));
 sky130_fd_sc_hd__xor2_2 _21360_ (.A(_03088_),
    .B(_03096_),
    .X(_03097_));
 sky130_fd_sc_hd__nand2_1 _21361_ (.A(_03009_),
    .B(_03054_),
    .Y(_03098_));
 sky130_fd_sc_hd__o21a_1 _21362_ (.A1(_03049_),
    .A2(_03055_),
    .B1(_03098_),
    .X(_03099_));
 sky130_fd_sc_hd__xnor2_2 _21363_ (.A(_03097_),
    .B(_03099_),
    .Y(_03100_));
 sky130_fd_sc_hd__xnor2_2 _21364_ (.A(_03083_),
    .B(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__nand2_1 _21365_ (.A(_03044_),
    .B(_03056_),
    .Y(_03102_));
 sky130_fd_sc_hd__o21a_1 _21366_ (.A1(_03043_),
    .A2(_03057_),
    .B1(_03102_),
    .X(_03103_));
 sky130_fd_sc_hd__xnor2_2 _21367_ (.A(_03101_),
    .B(_03103_),
    .Y(_03104_));
 sky130_fd_sc_hd__xor2_2 _21368_ (.A(_03074_),
    .B(_03104_),
    .X(_03105_));
 sky130_fd_sc_hd__or2b_1 _21369_ (.A(_03058_),
    .B_N(_03035_),
    .X(_03106_));
 sky130_fd_sc_hd__or2b_1 _21370_ (.A(_03059_),
    .B_N(_03034_),
    .X(_03107_));
 sky130_fd_sc_hd__and2_1 _21371_ (.A(_03106_),
    .B(_03107_),
    .X(_03108_));
 sky130_fd_sc_hd__xnor2_2 _21372_ (.A(_03105_),
    .B(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__and2b_1 _21373_ (.A_N(_03061_),
    .B(_03060_),
    .X(_03110_));
 sky130_fd_sc_hd__a21oi_2 _21374_ (.A1(_02897_),
    .A2(_03062_),
    .B1(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__xor2_2 _21375_ (.A(_03109_),
    .B(_03111_),
    .X(_03112_));
 sky130_fd_sc_hd__xor2_1 _21376_ (.A(_03072_),
    .B(_03112_),
    .X(_03113_));
 sky130_fd_sc_hd__or2_1 _21377_ (.A(net808),
    .B(_02638_),
    .X(_03114_));
 sky130_fd_sc_hd__o211a_1 _21378_ (.A1(_03070_),
    .A2(_03113_),
    .B1(_03114_),
    .C1(_02909_),
    .X(_00830_));
 sky130_fd_sc_hd__or2_1 _21379_ (.A(_03109_),
    .B(_03111_),
    .X(_03115_));
 sky130_fd_sc_hd__nand2_1 _21380_ (.A(_03072_),
    .B(_03112_),
    .Y(_03116_));
 sky130_fd_sc_hd__or2_2 _21381_ (.A(_03105_),
    .B(_03108_),
    .X(_03117_));
 sky130_fd_sc_hd__or2_1 _21382_ (.A(_03101_),
    .B(_03103_),
    .X(_03118_));
 sky130_fd_sc_hd__or2b_1 _21383_ (.A(_03104_),
    .B_N(_03074_),
    .X(_03119_));
 sky130_fd_sc_hd__or2b_1 _21384_ (.A(_03075_),
    .B_N(_03082_),
    .X(_03120_));
 sky130_fd_sc_hd__o21ai_1 _21385_ (.A1(_03076_),
    .A2(_03081_),
    .B1(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__clkbuf_4 _21386_ (.A(_03080_),
    .X(_03122_));
 sky130_fd_sc_hd__clkbuf_4 _21387_ (.A(_03077_),
    .X(_03123_));
 sky130_fd_sc_hd__a21o_1 _21388_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[8] ),
    .A2(_03122_),
    .B1(_03123_),
    .X(_03124_));
 sky130_fd_sc_hd__a21bo_1 _21389_ (.A1(_03084_),
    .A2(_03087_),
    .B1_N(_03085_),
    .X(_03125_));
 sky130_fd_sc_hd__nand2_1 _21390_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[9] ),
    .B(_03080_),
    .Y(_03126_));
 sky130_fd_sc_hd__or2_1 _21391_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[9] ),
    .B(_03080_),
    .X(_03127_));
 sky130_fd_sc_hd__nand2_1 _21392_ (.A(_03126_),
    .B(_03127_),
    .Y(_03128_));
 sky130_fd_sc_hd__xnor2_1 _21393_ (.A(_03125_),
    .B(_03128_),
    .Y(_03129_));
 sky130_fd_sc_hd__xor2_1 _21394_ (.A(_03124_),
    .B(_03129_),
    .X(_03130_));
 sky130_fd_sc_hd__a22o_1 _21395_ (.A1(\top_inst.grid_inst.data_path_wires[17][5] ),
    .A2(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[17][6] ),
    .X(_03131_));
 sky130_fd_sc_hd__and4_1 _21396_ (.A(\top_inst.grid_inst.data_path_wires[17][6] ),
    .B(\top_inst.grid_inst.data_path_wires[17][5] ),
    .C(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[3] ),
    .X(_03132_));
 sky130_fd_sc_hd__inv_2 _21397_ (.A(_03132_),
    .Y(_03133_));
 sky130_fd_sc_hd__and2_1 _21398_ (.A(_03131_),
    .B(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__nand2_4 _21399_ (.A(_02878_),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[2] ),
    .Y(_03135_));
 sky130_fd_sc_hd__xnor2_2 _21400_ (.A(_03134_),
    .B(_03135_),
    .Y(_03136_));
 sky130_fd_sc_hd__nand2_1 _21401_ (.A(\top_inst.grid_inst.data_path_wires[17][4] ),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[5] ),
    .Y(_03137_));
 sky130_fd_sc_hd__and2b_1 _21402_ (.A_N(\top_inst.grid_inst.data_path_wires[17][2] ),
    .B(_02897_),
    .X(_03138_));
 sky130_fd_sc_hd__nand2_1 _21403_ (.A(\top_inst.grid_inst.data_path_wires[17][3] ),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[6] ),
    .Y(_03139_));
 sky130_fd_sc_hd__xnor2_2 _21404_ (.A(_03138_),
    .B(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hd__xnor2_2 _21405_ (.A(_03137_),
    .B(_03140_),
    .Y(_03141_));
 sky130_fd_sc_hd__and3_1 _21406_ (.A(\top_inst.grid_inst.data_path_wires[17][2] ),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[6] ),
    .C(_03090_),
    .X(_03142_));
 sky130_fd_sc_hd__a31o_1 _21407_ (.A1(_02868_),
    .A2(_02893_),
    .A3(_03092_),
    .B1(_03142_),
    .X(_03143_));
 sky130_fd_sc_hd__xor2_2 _21408_ (.A(_03141_),
    .B(_03143_),
    .X(_03144_));
 sky130_fd_sc_hd__xnor2_2 _21409_ (.A(_03136_),
    .B(_03144_),
    .Y(_03145_));
 sky130_fd_sc_hd__and2_1 _21410_ (.A(_03093_),
    .B(_03095_),
    .X(_03146_));
 sky130_fd_sc_hd__a21o_1 _21411_ (.A1(_03088_),
    .A2(_03096_),
    .B1(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__xnor2_2 _21412_ (.A(_03145_),
    .B(_03147_),
    .Y(_03148_));
 sky130_fd_sc_hd__xnor2_1 _21413_ (.A(_03130_),
    .B(_03148_),
    .Y(_03149_));
 sky130_fd_sc_hd__and2b_1 _21414_ (.A_N(_03099_),
    .B(_03097_),
    .X(_03150_));
 sky130_fd_sc_hd__a21oi_1 _21415_ (.A1(_03083_),
    .A2(_03100_),
    .B1(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__xor2_1 _21416_ (.A(_03149_),
    .B(_03151_),
    .X(_03152_));
 sky130_fd_sc_hd__xnor2_1 _21417_ (.A(_03121_),
    .B(_03152_),
    .Y(_03153_));
 sky130_fd_sc_hd__a21oi_2 _21418_ (.A1(_03118_),
    .A2(_03119_),
    .B1(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__and3_1 _21419_ (.A(_03118_),
    .B(_03119_),
    .C(_03153_),
    .X(_03155_));
 sky130_fd_sc_hd__nor2_1 _21420_ (.A(_03154_),
    .B(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__xnor2_2 _21421_ (.A(_03117_),
    .B(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__a21oi_1 _21422_ (.A1(_03115_),
    .A2(_03116_),
    .B1(_03157_),
    .Y(_03158_));
 sky130_fd_sc_hd__a31o_1 _21423_ (.A1(_03115_),
    .A2(_03116_),
    .A3(_03157_),
    .B1(_01984_),
    .X(_03159_));
 sky130_fd_sc_hd__o221a_1 _21424_ (.A1(net924),
    .A2(_02491_),
    .B1(_03158_),
    .B2(_03159_),
    .C1(_02962_),
    .X(_00831_));
 sky130_fd_sc_hd__nor2_1 _21425_ (.A(_03149_),
    .B(_03151_),
    .Y(_03160_));
 sky130_fd_sc_hd__a21o_1 _21426_ (.A1(_03121_),
    .A2(_03152_),
    .B1(_03160_),
    .X(_03161_));
 sky130_fd_sc_hd__a32o_1 _21427_ (.A1(_03125_),
    .A2(_03126_),
    .A3(_03127_),
    .B1(_03129_),
    .B2(_03124_),
    .X(_03162_));
 sky130_fd_sc_hd__a21o_1 _21428_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[9] ),
    .A2(_03122_),
    .B1(_03123_),
    .X(_03163_));
 sky130_fd_sc_hd__a31o_1 _21429_ (.A1(_02878_),
    .A2(_02887_),
    .A3(_03131_),
    .B1(_03132_),
    .X(_03164_));
 sky130_fd_sc_hd__xnor2_2 _21430_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[10] ),
    .B(_03080_),
    .Y(_03165_));
 sky130_fd_sc_hd__xnor2_2 _21431_ (.A(_03164_),
    .B(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__xnor2_2 _21432_ (.A(_03163_),
    .B(_03166_),
    .Y(_03167_));
 sky130_fd_sc_hd__and3_1 _21433_ (.A(\top_inst.grid_inst.data_path_wires[17][7] ),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[4] ),
    .C(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[3] ),
    .X(_03168_));
 sky130_fd_sc_hd__a22o_1 _21434_ (.A1(\top_inst.grid_inst.data_path_wires[17][6] ),
    .A2(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[17][7] ),
    .X(_03169_));
 sky130_fd_sc_hd__a21bo_1 _21435_ (.A1(_02875_),
    .A2(_03168_),
    .B1_N(_03169_),
    .X(_03170_));
 sky130_fd_sc_hd__xor2_2 _21436_ (.A(_03135_),
    .B(_03170_),
    .X(_03171_));
 sky130_fd_sc_hd__nand2_1 _21437_ (.A(_02873_),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[5] ),
    .Y(_03172_));
 sky130_fd_sc_hd__and2b_1 _21438_ (.A_N(\top_inst.grid_inst.data_path_wires[17][3] ),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[7] ),
    .X(_03173_));
 sky130_fd_sc_hd__nand2_1 _21439_ (.A(\top_inst.grid_inst.data_path_wires[17][4] ),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[6] ),
    .Y(_03174_));
 sky130_fd_sc_hd__xnor2_2 _21440_ (.A(_03173_),
    .B(_03174_),
    .Y(_03175_));
 sky130_fd_sc_hd__xnor2_2 _21441_ (.A(_03172_),
    .B(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__and3_1 _21442_ (.A(\top_inst.grid_inst.data_path_wires[17][3] ),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[6] ),
    .C(_03138_),
    .X(_03177_));
 sky130_fd_sc_hd__a31o_1 _21443_ (.A1(_02871_),
    .A2(_02893_),
    .A3(_03140_),
    .B1(_03177_),
    .X(_03178_));
 sky130_fd_sc_hd__xor2_2 _21444_ (.A(_03176_),
    .B(_03178_),
    .X(_03179_));
 sky130_fd_sc_hd__xnor2_2 _21445_ (.A(_03171_),
    .B(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__nand2_1 _21446_ (.A(_03141_),
    .B(_03143_),
    .Y(_03181_));
 sky130_fd_sc_hd__a21boi_2 _21447_ (.A1(_03136_),
    .A2(_03144_),
    .B1_N(_03181_),
    .Y(_03182_));
 sky130_fd_sc_hd__xnor2_2 _21448_ (.A(_03180_),
    .B(_03182_),
    .Y(_03183_));
 sky130_fd_sc_hd__xnor2_2 _21449_ (.A(_03167_),
    .B(_03183_),
    .Y(_03184_));
 sky130_fd_sc_hd__and2b_1 _21450_ (.A_N(_03145_),
    .B(_03147_),
    .X(_03185_));
 sky130_fd_sc_hd__a21oi_2 _21451_ (.A1(_03130_),
    .A2(_03148_),
    .B1(_03185_),
    .Y(_03186_));
 sky130_fd_sc_hd__xor2_2 _21452_ (.A(_03184_),
    .B(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__xnor2_2 _21453_ (.A(_03162_),
    .B(_03187_),
    .Y(_03188_));
 sky130_fd_sc_hd__xnor2_2 _21454_ (.A(_03161_),
    .B(_03188_),
    .Y(_03189_));
 sky130_fd_sc_hd__xor2_2 _21455_ (.A(_03154_),
    .B(_03189_),
    .X(_03190_));
 sky130_fd_sc_hd__a21boi_2 _21456_ (.A1(_03117_),
    .A2(_03115_),
    .B1_N(_03156_),
    .Y(_03191_));
 sky130_fd_sc_hd__a31o_1 _21457_ (.A1(_03072_),
    .A2(_03112_),
    .A3(_03157_),
    .B1(_03191_),
    .X(_03192_));
 sky130_fd_sc_hd__nand2_1 _21458_ (.A(_03190_),
    .B(_03192_),
    .Y(_03193_));
 sky130_fd_sc_hd__o21a_1 _21459_ (.A1(_03190_),
    .A2(_03192_),
    .B1(_10831_),
    .X(_03194_));
 sky130_fd_sc_hd__a22o_1 _21460_ (.A1(\top_inst.deskew_buff_inst.col_input[74] ),
    .A2(_05731_),
    .B1(_03193_),
    .B2(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__and2_1 _21461_ (.A(_02135_),
    .B(_03195_),
    .X(_03196_));
 sky130_fd_sc_hd__clkbuf_1 _21462_ (.A(_03196_),
    .X(_00832_));
 sky130_fd_sc_hd__nand2_1 _21463_ (.A(_03154_),
    .B(_03189_),
    .Y(_03197_));
 sky130_fd_sc_hd__or2b_1 _21464_ (.A(_03188_),
    .B_N(_03161_),
    .X(_03198_));
 sky130_fd_sc_hd__or2b_1 _21465_ (.A(_03165_),
    .B_N(_03164_),
    .X(_03199_));
 sky130_fd_sc_hd__a21bo_1 _21466_ (.A1(_03163_),
    .A2(_03166_),
    .B1_N(_03199_),
    .X(_03200_));
 sky130_fd_sc_hd__a21o_1 _21467_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[10] ),
    .A2(_03080_),
    .B1(_03123_),
    .X(_03201_));
 sky130_fd_sc_hd__a32o_1 _21468_ (.A1(_02878_),
    .A2(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[2] ),
    .A3(_03169_),
    .B1(_03168_),
    .B2(_02875_),
    .X(_03202_));
 sky130_fd_sc_hd__xnor2_1 _21469_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[11] ),
    .B(_03079_),
    .Y(_03203_));
 sky130_fd_sc_hd__xnor2_1 _21470_ (.A(_03202_),
    .B(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__and2_1 _21471_ (.A(_03201_),
    .B(_03204_),
    .X(_03205_));
 sky130_fd_sc_hd__nor2_1 _21472_ (.A(_03201_),
    .B(_03204_),
    .Y(_03206_));
 sky130_fd_sc_hd__or2_1 _21473_ (.A(_03205_),
    .B(_03206_),
    .X(_03207_));
 sky130_fd_sc_hd__o21ai_1 _21474_ (.A1(_02891_),
    .A2(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[3] ),
    .B1(_02878_),
    .Y(_03208_));
 sky130_fd_sc_hd__nor2_2 _21475_ (.A(_03168_),
    .B(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__xnor2_4 _21476_ (.A(_03135_),
    .B(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__nand2_1 _21477_ (.A(\top_inst.grid_inst.data_path_wires[17][6] ),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[5] ),
    .Y(_03211_));
 sky130_fd_sc_hd__and2b_1 _21478_ (.A_N(\top_inst.grid_inst.data_path_wires[17][4] ),
    .B(_02897_),
    .X(_03212_));
 sky130_fd_sc_hd__nand2_1 _21479_ (.A(\top_inst.grid_inst.data_path_wires[17][5] ),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[6] ),
    .Y(_03213_));
 sky130_fd_sc_hd__xnor2_2 _21480_ (.A(_03212_),
    .B(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__xnor2_2 _21481_ (.A(_03211_),
    .B(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__and3_1 _21482_ (.A(\top_inst.grid_inst.data_path_wires[17][4] ),
    .B(_02895_),
    .C(_03173_),
    .X(_03216_));
 sky130_fd_sc_hd__a31o_1 _21483_ (.A1(_02873_),
    .A2(_02893_),
    .A3(_03175_),
    .B1(_03216_),
    .X(_03217_));
 sky130_fd_sc_hd__xor2_2 _21484_ (.A(_03215_),
    .B(_03217_),
    .X(_03218_));
 sky130_fd_sc_hd__xnor2_2 _21485_ (.A(_03210_),
    .B(_03218_),
    .Y(_03219_));
 sky130_fd_sc_hd__and2_1 _21486_ (.A(_03176_),
    .B(_03178_),
    .X(_03220_));
 sky130_fd_sc_hd__a21oi_2 _21487_ (.A1(_03171_),
    .A2(_03179_),
    .B1(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__xnor2_2 _21488_ (.A(_03219_),
    .B(_03221_),
    .Y(_03222_));
 sky130_fd_sc_hd__xor2_2 _21489_ (.A(_03207_),
    .B(_03222_),
    .X(_03223_));
 sky130_fd_sc_hd__or2_1 _21490_ (.A(_03180_),
    .B(_03182_),
    .X(_03224_));
 sky130_fd_sc_hd__o21a_1 _21491_ (.A1(_03167_),
    .A2(_03183_),
    .B1(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__xor2_2 _21492_ (.A(_03223_),
    .B(_03225_),
    .X(_03226_));
 sky130_fd_sc_hd__xor2_2 _21493_ (.A(_03200_),
    .B(_03226_),
    .X(_03227_));
 sky130_fd_sc_hd__nor2_1 _21494_ (.A(_03184_),
    .B(_03186_),
    .Y(_03228_));
 sky130_fd_sc_hd__a21oi_2 _21495_ (.A1(_03162_),
    .A2(_03187_),
    .B1(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__xor2_2 _21496_ (.A(_03227_),
    .B(_03229_),
    .X(_03230_));
 sky130_fd_sc_hd__xnor2_2 _21497_ (.A(_03198_),
    .B(_03230_),
    .Y(_03231_));
 sky130_fd_sc_hd__a21oi_1 _21498_ (.A1(_03197_),
    .A2(_03193_),
    .B1(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__and3_1 _21499_ (.A(_03197_),
    .B(_03193_),
    .C(_03231_),
    .X(_03233_));
 sky130_fd_sc_hd__or2_1 _21500_ (.A(net753),
    .B(_05316_),
    .X(_03234_));
 sky130_fd_sc_hd__o311a_1 _21501_ (.A1(_09787_),
    .A2(_03232_),
    .A3(_03233_),
    .B1(_03234_),
    .C1(_09806_),
    .X(_00833_));
 sky130_fd_sc_hd__and2_1 _21502_ (.A(_03190_),
    .B(_03231_),
    .X(_03235_));
 sky130_fd_sc_hd__and3_1 _21503_ (.A(_03112_),
    .B(_03157_),
    .C(_03235_),
    .X(_03236_));
 sky130_fd_sc_hd__a21boi_2 _21504_ (.A1(_03198_),
    .A2(_03197_),
    .B1_N(_03230_),
    .Y(_03237_));
 sky130_fd_sc_hd__a221oi_4 _21505_ (.A1(_03191_),
    .A2(_03235_),
    .B1(_03236_),
    .B2(_03072_),
    .C1(_03237_),
    .Y(_03238_));
 sky130_fd_sc_hd__nor2_1 _21506_ (.A(_03227_),
    .B(_03229_),
    .Y(_03239_));
 sky130_fd_sc_hd__or2b_1 _21507_ (.A(_03225_),
    .B_N(_03223_),
    .X(_03240_));
 sky130_fd_sc_hd__or2b_1 _21508_ (.A(_03226_),
    .B_N(_03200_),
    .X(_03241_));
 sky130_fd_sc_hd__or2b_1 _21509_ (.A(_03203_),
    .B_N(_03202_),
    .X(_03242_));
 sky130_fd_sc_hd__a21bo_1 _21510_ (.A1(_03201_),
    .A2(_03204_),
    .B1_N(_03242_),
    .X(_03243_));
 sky130_fd_sc_hd__a21o_1 _21511_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[11] ),
    .A2(_03122_),
    .B1(_03123_),
    .X(_03244_));
 sky130_fd_sc_hd__o21ba_1 _21512_ (.A1(_03135_),
    .A2(_03208_),
    .B1_N(_03168_),
    .X(_03245_));
 sky130_fd_sc_hd__clkbuf_4 _21513_ (.A(_03245_),
    .X(_03246_));
 sky130_fd_sc_hd__xnor2_1 _21514_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[12] ),
    .B(_03080_),
    .Y(_03247_));
 sky130_fd_sc_hd__xor2_1 _21515_ (.A(_03246_),
    .B(_03247_),
    .X(_03248_));
 sky130_fd_sc_hd__and2_1 _21516_ (.A(_03244_),
    .B(_03248_),
    .X(_03249_));
 sky130_fd_sc_hd__nor2_1 _21517_ (.A(_03244_),
    .B(_03248_),
    .Y(_03250_));
 sky130_fd_sc_hd__or2_1 _21518_ (.A(_03249_),
    .B(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__and2_1 _21519_ (.A(\top_inst.grid_inst.data_path_wires[17][7] ),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[5] ),
    .X(_03252_));
 sky130_fd_sc_hd__buf_2 _21520_ (.A(_03252_),
    .X(_03253_));
 sky130_fd_sc_hd__and2b_1 _21521_ (.A_N(\top_inst.grid_inst.data_path_wires[17][5] ),
    .B(_02897_),
    .X(_03254_));
 sky130_fd_sc_hd__nand2_1 _21522_ (.A(\top_inst.grid_inst.data_path_wires[17][6] ),
    .B(_02895_),
    .Y(_03255_));
 sky130_fd_sc_hd__xor2_1 _21523_ (.A(_03254_),
    .B(_03255_),
    .X(_03256_));
 sky130_fd_sc_hd__xnor2_2 _21524_ (.A(_03253_),
    .B(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__and3_1 _21525_ (.A(_02873_),
    .B(_02895_),
    .C(_03212_),
    .X(_03258_));
 sky130_fd_sc_hd__a31o_1 _21526_ (.A1(_02875_),
    .A2(_02893_),
    .A3(_03214_),
    .B1(_03258_),
    .X(_03259_));
 sky130_fd_sc_hd__xor2_2 _21527_ (.A(_03257_),
    .B(_03259_),
    .X(_03260_));
 sky130_fd_sc_hd__xnor2_1 _21528_ (.A(_03210_),
    .B(_03260_),
    .Y(_03261_));
 sky130_fd_sc_hd__and2_1 _21529_ (.A(_03215_),
    .B(_03217_),
    .X(_03262_));
 sky130_fd_sc_hd__a21oi_1 _21530_ (.A1(_03210_),
    .A2(_03218_),
    .B1(_03262_),
    .Y(_03263_));
 sky130_fd_sc_hd__xnor2_1 _21531_ (.A(_03261_),
    .B(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hd__xor2_1 _21532_ (.A(_03251_),
    .B(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__o32a_1 _21533_ (.A1(_03205_),
    .A2(_03206_),
    .A3(_03222_),
    .B1(_03221_),
    .B2(_03219_),
    .X(_03266_));
 sky130_fd_sc_hd__xnor2_1 _21534_ (.A(_03265_),
    .B(_03266_),
    .Y(_03267_));
 sky130_fd_sc_hd__xnor2_1 _21535_ (.A(_03243_),
    .B(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__a21o_1 _21536_ (.A1(_03240_),
    .A2(_03241_),
    .B1(_03268_),
    .X(_03269_));
 sky130_fd_sc_hd__nand3_1 _21537_ (.A(_03240_),
    .B(_03241_),
    .C(_03268_),
    .Y(_03270_));
 sky130_fd_sc_hd__and2_1 _21538_ (.A(_03269_),
    .B(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__xor2_2 _21539_ (.A(_03239_),
    .B(_03271_),
    .X(_03272_));
 sky130_fd_sc_hd__xnor2_1 _21540_ (.A(_03238_),
    .B(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__or2_1 _21541_ (.A(net839),
    .B(_02638_),
    .X(_03274_));
 sky130_fd_sc_hd__o211a_1 _21542_ (.A1(_03070_),
    .A2(_03273_),
    .B1(_03274_),
    .C1(_02909_),
    .X(_00834_));
 sky130_fd_sc_hd__a31o_1 _21543_ (.A1(_03190_),
    .A2(_03192_),
    .A3(_03231_),
    .B1(_03237_),
    .X(_03275_));
 sky130_fd_sc_hd__nand2_1 _21544_ (.A(_03239_),
    .B(_03271_),
    .Y(_03276_));
 sky130_fd_sc_hd__a21bo_1 _21545_ (.A1(_03275_),
    .A2(_03272_),
    .B1_N(_03276_),
    .X(_03277_));
 sky130_fd_sc_hd__buf_2 _21546_ (.A(_03246_),
    .X(_03278_));
 sky130_fd_sc_hd__clkbuf_4 _21547_ (.A(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__o21bai_1 _21548_ (.A1(_03279_),
    .A2(_03247_),
    .B1_N(_03249_),
    .Y(_03280_));
 sky130_fd_sc_hd__a21o_1 _21549_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[12] ),
    .A2(_03122_),
    .B1(_03123_),
    .X(_03281_));
 sky130_fd_sc_hd__xnor2_1 _21550_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[13] ),
    .B(_03080_),
    .Y(_03282_));
 sky130_fd_sc_hd__xor2_1 _21551_ (.A(_03245_),
    .B(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__and2_1 _21552_ (.A(_03281_),
    .B(_03283_),
    .X(_03284_));
 sky130_fd_sc_hd__nor2_1 _21553_ (.A(_03281_),
    .B(_03283_),
    .Y(_03285_));
 sky130_fd_sc_hd__or2_1 _21554_ (.A(_03284_),
    .B(_03285_),
    .X(_03286_));
 sky130_fd_sc_hd__nand2_1 _21555_ (.A(\top_inst.grid_inst.data_path_wires[17][7] ),
    .B(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[6] ),
    .Y(_03287_));
 sky130_fd_sc_hd__nand2b_1 _21556_ (.A_N(\top_inst.grid_inst.data_path_wires[17][6] ),
    .B(_02897_),
    .Y(_03288_));
 sky130_fd_sc_hd__xnor2_1 _21557_ (.A(_03287_),
    .B(_03288_),
    .Y(_03289_));
 sky130_fd_sc_hd__xnor2_2 _21558_ (.A(_03253_),
    .B(_03289_),
    .Y(_03290_));
 sky130_fd_sc_hd__or2b_1 _21559_ (.A(_03254_),
    .B_N(_03255_),
    .X(_03291_));
 sky130_fd_sc_hd__and3_1 _21560_ (.A(_02875_),
    .B(_02895_),
    .C(_03254_),
    .X(_03292_));
 sky130_fd_sc_hd__a21o_1 _21561_ (.A1(_03253_),
    .A2(_03291_),
    .B1(_03292_),
    .X(_03293_));
 sky130_fd_sc_hd__xor2_2 _21562_ (.A(_03290_),
    .B(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__xnor2_2 _21563_ (.A(_03210_),
    .B(_03294_),
    .Y(_03295_));
 sky130_fd_sc_hd__and2_1 _21564_ (.A(_03257_),
    .B(_03259_),
    .X(_03296_));
 sky130_fd_sc_hd__a21oi_2 _21565_ (.A1(_03210_),
    .A2(_03260_),
    .B1(_03296_),
    .Y(_03297_));
 sky130_fd_sc_hd__xnor2_2 _21566_ (.A(_03295_),
    .B(_03297_),
    .Y(_03298_));
 sky130_fd_sc_hd__xor2_2 _21567_ (.A(_03286_),
    .B(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__o32a_1 _21568_ (.A1(_03249_),
    .A2(_03250_),
    .A3(_03264_),
    .B1(_03263_),
    .B2(_03261_),
    .X(_03300_));
 sky130_fd_sc_hd__xor2_1 _21569_ (.A(_03299_),
    .B(_03300_),
    .X(_03301_));
 sky130_fd_sc_hd__xor2_1 _21570_ (.A(_03280_),
    .B(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__and2b_1 _21571_ (.A_N(_03266_),
    .B(_03265_),
    .X(_03303_));
 sky130_fd_sc_hd__a21oi_1 _21572_ (.A1(_03243_),
    .A2(_03267_),
    .B1(_03303_),
    .Y(_03304_));
 sky130_fd_sc_hd__nor2_1 _21573_ (.A(_03302_),
    .B(_03304_),
    .Y(_03305_));
 sky130_fd_sc_hd__and2_1 _21574_ (.A(_03302_),
    .B(_03304_),
    .X(_03306_));
 sky130_fd_sc_hd__nor2_1 _21575_ (.A(_03305_),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__xnor2_1 _21576_ (.A(_03269_),
    .B(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hd__xor2_1 _21577_ (.A(_03277_),
    .B(_03308_),
    .X(_03309_));
 sky130_fd_sc_hd__or2_1 _21578_ (.A(net818),
    .B(_02638_),
    .X(_03310_));
 sky130_fd_sc_hd__o211a_1 _21579_ (.A1(_03070_),
    .A2(_03309_),
    .B1(_03310_),
    .C1(_02909_),
    .X(_00835_));
 sky130_fd_sc_hd__clkbuf_4 _21580_ (.A(_04873_),
    .X(_03311_));
 sky130_fd_sc_hd__or2b_1 _21581_ (.A(_03300_),
    .B_N(_03299_),
    .X(_03312_));
 sky130_fd_sc_hd__or2b_1 _21582_ (.A(_03301_),
    .B_N(_03280_),
    .X(_03313_));
 sky130_fd_sc_hd__o21bai_2 _21583_ (.A1(_03279_),
    .A2(_03282_),
    .B1_N(_03284_),
    .Y(_03314_));
 sky130_fd_sc_hd__a21o_1 _21584_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[13] ),
    .A2(_03122_),
    .B1(_03123_),
    .X(_03315_));
 sky130_fd_sc_hd__xnor2_1 _21585_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[14] ),
    .B(_03080_),
    .Y(_03316_));
 sky130_fd_sc_hd__nor2_1 _21586_ (.A(_03246_),
    .B(_03316_),
    .Y(_03317_));
 sky130_fd_sc_hd__and2_1 _21587_ (.A(_03246_),
    .B(_03316_),
    .X(_03318_));
 sky130_fd_sc_hd__nor2_1 _21588_ (.A(_03317_),
    .B(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__xnor2_2 _21589_ (.A(_03315_),
    .B(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__and2_1 _21590_ (.A(_03290_),
    .B(_03293_),
    .X(_03321_));
 sky130_fd_sc_hd__a21oi_2 _21591_ (.A1(_03210_),
    .A2(_03294_),
    .B1(_03321_),
    .Y(_03322_));
 sky130_fd_sc_hd__nand2_1 _21592_ (.A(_03287_),
    .B(_03288_),
    .Y(_03323_));
 sky130_fd_sc_hd__nor2_1 _21593_ (.A(_03287_),
    .B(_03288_),
    .Y(_03324_));
 sky130_fd_sc_hd__a21o_1 _21594_ (.A1(_03253_),
    .A2(_03323_),
    .B1(_03324_),
    .X(_03325_));
 sky130_fd_sc_hd__nand2_1 _21595_ (.A(_02895_),
    .B(_03253_),
    .Y(_03326_));
 sky130_fd_sc_hd__mux2_1 _21596_ (.A0(_02897_),
    .A1(_02895_),
    .S(_02878_),
    .X(_03327_));
 sky130_fd_sc_hd__nor2_1 _21597_ (.A(_03253_),
    .B(_03327_),
    .Y(_03328_));
 sky130_fd_sc_hd__a21oi_2 _21598_ (.A1(_03325_),
    .A2(_03326_),
    .B1(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__xnor2_2 _21599_ (.A(_03210_),
    .B(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__xor2_2 _21600_ (.A(_03322_),
    .B(_03330_),
    .X(_03331_));
 sky130_fd_sc_hd__xnor2_2 _21601_ (.A(_03320_),
    .B(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__o32a_1 _21602_ (.A1(_03284_),
    .A2(_03285_),
    .A3(_03298_),
    .B1(_03297_),
    .B2(_03295_),
    .X(_03333_));
 sky130_fd_sc_hd__xnor2_2 _21603_ (.A(_03332_),
    .B(_03333_),
    .Y(_03334_));
 sky130_fd_sc_hd__xnor2_1 _21604_ (.A(_03314_),
    .B(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__a21o_1 _21605_ (.A1(_03312_),
    .A2(_03313_),
    .B1(_03335_),
    .X(_03336_));
 sky130_fd_sc_hd__nand3_1 _21606_ (.A(_03312_),
    .B(_03313_),
    .C(_03335_),
    .Y(_03337_));
 sky130_fd_sc_hd__and2_1 _21607_ (.A(_03336_),
    .B(_03337_),
    .X(_03338_));
 sky130_fd_sc_hd__xor2_1 _21608_ (.A(_03305_),
    .B(_03338_),
    .X(_03339_));
 sky130_fd_sc_hd__and2_1 _21609_ (.A(_03272_),
    .B(_03308_),
    .X(_03340_));
 sky130_fd_sc_hd__a21boi_1 _21610_ (.A1(_03269_),
    .A2(_03276_),
    .B1_N(_03307_),
    .Y(_03341_));
 sky130_fd_sc_hd__a21o_1 _21611_ (.A1(_03275_),
    .A2(_03340_),
    .B1(_03341_),
    .X(_03342_));
 sky130_fd_sc_hd__nand2_1 _21612_ (.A(_03339_),
    .B(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__o21a_1 _21613_ (.A1(_03339_),
    .A2(_03342_),
    .B1(_10831_),
    .X(_03344_));
 sky130_fd_sc_hd__a22o_1 _21614_ (.A1(\top_inst.deskew_buff_inst.col_input[78] ),
    .A2(_05731_),
    .B1(_03343_),
    .B2(_03344_),
    .X(_03345_));
 sky130_fd_sc_hd__and2_1 _21615_ (.A(_03311_),
    .B(_03345_),
    .X(_03346_));
 sky130_fd_sc_hd__clkbuf_1 _21616_ (.A(_03346_),
    .X(_00836_));
 sky130_fd_sc_hd__nand2_1 _21617_ (.A(_03305_),
    .B(_03338_),
    .Y(_03347_));
 sky130_fd_sc_hd__a21o_1 _21618_ (.A1(_03315_),
    .A2(_03319_),
    .B1(_03317_),
    .X(_03348_));
 sky130_fd_sc_hd__nor2_1 _21619_ (.A(_03322_),
    .B(_03330_),
    .Y(_03349_));
 sky130_fd_sc_hd__and2b_1 _21620_ (.A_N(_03320_),
    .B(_03331_),
    .X(_03350_));
 sky130_fd_sc_hd__nor2_1 _21621_ (.A(_03210_),
    .B(_03329_),
    .Y(_03351_));
 sky130_fd_sc_hd__a21o_1 _21622_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[14] ),
    .A2(_03122_),
    .B1(_03123_),
    .X(_03352_));
 sky130_fd_sc_hd__xnor2_1 _21623_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[15] ),
    .B(_03080_),
    .Y(_03353_));
 sky130_fd_sc_hd__xor2_1 _21624_ (.A(_03245_),
    .B(_03353_),
    .X(_03354_));
 sky130_fd_sc_hd__xnor2_1 _21625_ (.A(_03352_),
    .B(_03354_),
    .Y(_03355_));
 sky130_fd_sc_hd__or2_1 _21626_ (.A(_03351_),
    .B(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__nand2_1 _21627_ (.A(_03351_),
    .B(_03355_),
    .Y(_03357_));
 sky130_fd_sc_hd__and2_1 _21628_ (.A(_03356_),
    .B(_03357_),
    .X(_03358_));
 sky130_fd_sc_hd__o21a_1 _21629_ (.A1(_03349_),
    .A2(_03350_),
    .B1(_03358_),
    .X(_03359_));
 sky130_fd_sc_hd__or3_1 _21630_ (.A(_03349_),
    .B(_03350_),
    .C(_03358_),
    .X(_03360_));
 sky130_fd_sc_hd__and2b_1 _21631_ (.A_N(_03359_),
    .B(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__xnor2_2 _21632_ (.A(_03348_),
    .B(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__and2b_1 _21633_ (.A_N(_03333_),
    .B(_03332_),
    .X(_03363_));
 sky130_fd_sc_hd__a21oi_2 _21634_ (.A1(_03314_),
    .A2(_03334_),
    .B1(_03363_),
    .Y(_03364_));
 sky130_fd_sc_hd__xor2_2 _21635_ (.A(_03362_),
    .B(_03364_),
    .X(_03365_));
 sky130_fd_sc_hd__xnor2_1 _21636_ (.A(_03336_),
    .B(_03365_),
    .Y(_03366_));
 sky130_fd_sc_hd__a21oi_1 _21637_ (.A1(_03347_),
    .A2(_03343_),
    .B1(_03366_),
    .Y(_03367_));
 sky130_fd_sc_hd__and3_1 _21638_ (.A(_03347_),
    .B(_03343_),
    .C(_03366_),
    .X(_03368_));
 sky130_fd_sc_hd__or2_1 _21639_ (.A(net544),
    .B(_05316_),
    .X(_03369_));
 sky130_fd_sc_hd__o311a_1 _21640_ (.A1(_09787_),
    .A2(_03367_),
    .A3(_03368_),
    .B1(_03369_),
    .C1(_09806_),
    .X(_00837_));
 sky130_fd_sc_hd__nor2_1 _21641_ (.A(_03362_),
    .B(_03364_),
    .Y(_03370_));
 sky130_fd_sc_hd__nor2_1 _21642_ (.A(_03279_),
    .B(_03353_),
    .Y(_03371_));
 sky130_fd_sc_hd__a21o_1 _21643_ (.A1(_03352_),
    .A2(_03354_),
    .B1(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__nand3b_1 _21644_ (.A_N(_03210_),
    .B(_03325_),
    .C(_03326_),
    .Y(_03373_));
 sky130_fd_sc_hd__and2b_1 _21645_ (.A_N(_03210_),
    .B(_03328_),
    .X(_03374_));
 sky130_fd_sc_hd__buf_2 _21646_ (.A(_03374_),
    .X(_03375_));
 sky130_fd_sc_hd__buf_4 _21647_ (.A(_03122_),
    .X(_03376_));
 sky130_fd_sc_hd__a21o_1 _21648_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[15] ),
    .A2(_03376_),
    .B1(_03123_),
    .X(_03377_));
 sky130_fd_sc_hd__xnor2_1 _21649_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[16] ),
    .B(_03122_),
    .Y(_03378_));
 sky130_fd_sc_hd__nor2_1 _21650_ (.A(_03246_),
    .B(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__and2_1 _21651_ (.A(_03246_),
    .B(_03378_),
    .X(_03380_));
 sky130_fd_sc_hd__nor2_1 _21652_ (.A(_03379_),
    .B(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__xnor2_1 _21653_ (.A(_03377_),
    .B(_03381_),
    .Y(_03382_));
 sky130_fd_sc_hd__xnor2_1 _21654_ (.A(_03375_),
    .B(_03382_),
    .Y(_03383_));
 sky130_fd_sc_hd__a21oi_1 _21655_ (.A1(_03356_),
    .A2(_03373_),
    .B1(_03383_),
    .Y(_03384_));
 sky130_fd_sc_hd__and3_1 _21656_ (.A(_03356_),
    .B(_03373_),
    .C(_03383_),
    .X(_03385_));
 sky130_fd_sc_hd__nor2_1 _21657_ (.A(_03384_),
    .B(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__xnor2_1 _21658_ (.A(_03372_),
    .B(_03386_),
    .Y(_03387_));
 sky130_fd_sc_hd__a21oi_1 _21659_ (.A1(_03348_),
    .A2(_03360_),
    .B1(_03359_),
    .Y(_03388_));
 sky130_fd_sc_hd__or2_2 _21660_ (.A(_03387_),
    .B(_03388_),
    .X(_03389_));
 sky130_fd_sc_hd__nand2_1 _21661_ (.A(_03387_),
    .B(_03388_),
    .Y(_03390_));
 sky130_fd_sc_hd__and2_1 _21662_ (.A(_03389_),
    .B(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__nand2_1 _21663_ (.A(_03370_),
    .B(_03391_),
    .Y(_03392_));
 sky130_fd_sc_hd__or2_1 _21664_ (.A(_03370_),
    .B(_03391_),
    .X(_03393_));
 sky130_fd_sc_hd__nand2_1 _21665_ (.A(_03392_),
    .B(_03393_),
    .Y(_03394_));
 sky130_fd_sc_hd__and2_1 _21666_ (.A(_03339_),
    .B(_03366_),
    .X(_03395_));
 sky130_fd_sc_hd__nand2_1 _21667_ (.A(_03340_),
    .B(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__nand2_1 _21668_ (.A(_03341_),
    .B(_03395_),
    .Y(_03397_));
 sky130_fd_sc_hd__a21bo_1 _21669_ (.A1(_03336_),
    .A2(_03347_),
    .B1_N(_03365_),
    .X(_03398_));
 sky130_fd_sc_hd__o211a_2 _21670_ (.A1(_03238_),
    .A2(_03396_),
    .B1(_03397_),
    .C1(_03398_),
    .X(_03399_));
 sky130_fd_sc_hd__xor2_1 _21671_ (.A(_03394_),
    .B(_03399_),
    .X(_03400_));
 sky130_fd_sc_hd__or2_1 _21672_ (.A(net411),
    .B(_02638_),
    .X(_03401_));
 sky130_fd_sc_hd__o211a_1 _21673_ (.A1(_03070_),
    .A2(_03400_),
    .B1(_03401_),
    .C1(_02909_),
    .X(_00838_));
 sky130_fd_sc_hd__o21a_1 _21674_ (.A1(_03394_),
    .A2(_03399_),
    .B1(_03392_),
    .X(_03402_));
 sky130_fd_sc_hd__a21o_1 _21675_ (.A1(_03377_),
    .A2(_03381_),
    .B1(_03379_),
    .X(_03403_));
 sky130_fd_sc_hd__or2b_1 _21676_ (.A(_03375_),
    .B_N(_03382_),
    .X(_03404_));
 sky130_fd_sc_hd__a21oi_2 _21677_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[16] ),
    .A2(_03376_),
    .B1(_03123_),
    .Y(_03405_));
 sky130_fd_sc_hd__xnor2_1 _21678_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[17] ),
    .B(_03122_),
    .Y(_03406_));
 sky130_fd_sc_hd__nor2_1 _21679_ (.A(_03246_),
    .B(_03406_),
    .Y(_03407_));
 sky130_fd_sc_hd__and2_1 _21680_ (.A(_03246_),
    .B(_03406_),
    .X(_03408_));
 sky130_fd_sc_hd__nor2_1 _21681_ (.A(_03407_),
    .B(_03408_),
    .Y(_03409_));
 sky130_fd_sc_hd__xnor2_2 _21682_ (.A(_03405_),
    .B(_03409_),
    .Y(_03410_));
 sky130_fd_sc_hd__xnor2_1 _21683_ (.A(_03404_),
    .B(_03410_),
    .Y(_03411_));
 sky130_fd_sc_hd__xnor2_1 _21684_ (.A(_03403_),
    .B(_03411_),
    .Y(_03412_));
 sky130_fd_sc_hd__a21oi_1 _21685_ (.A1(_03372_),
    .A2(_03386_),
    .B1(_03384_),
    .Y(_03413_));
 sky130_fd_sc_hd__nor2_1 _21686_ (.A(_03412_),
    .B(_03413_),
    .Y(_03414_));
 sky130_fd_sc_hd__nand2_1 _21687_ (.A(_03412_),
    .B(_03413_),
    .Y(_03415_));
 sky130_fd_sc_hd__or2b_1 _21688_ (.A(_03414_),
    .B_N(_03415_),
    .X(_03416_));
 sky130_fd_sc_hd__xor2_2 _21689_ (.A(_03389_),
    .B(_03416_),
    .X(_03417_));
 sky130_fd_sc_hd__nor2_1 _21690_ (.A(_03402_),
    .B(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__a2111o_1 _21691_ (.A1(_03402_),
    .A2(_03417_),
    .B1(_03418_),
    .C1(_05309_),
    .D1(_04861_),
    .X(_03419_));
 sky130_fd_sc_hd__o211a_1 _21692_ (.A1(net891),
    .A2(_06169_),
    .B1(_03419_),
    .C1(_02909_),
    .X(_00839_));
 sky130_fd_sc_hd__o21bai_2 _21693_ (.A1(_03405_),
    .A2(_03408_),
    .B1_N(_03407_),
    .Y(_03420_));
 sky130_fd_sc_hd__buf_4 _21694_ (.A(_03376_),
    .X(_03421_));
 sky130_fd_sc_hd__buf_4 _21695_ (.A(_03123_),
    .X(_03422_));
 sky130_fd_sc_hd__a21oi_2 _21696_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[17] ),
    .A2(_03421_),
    .B1(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__xnor2_1 _21697_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[18] ),
    .B(_03376_),
    .Y(_03424_));
 sky130_fd_sc_hd__nor2_1 _21698_ (.A(_03279_),
    .B(_03424_),
    .Y(_03425_));
 sky130_fd_sc_hd__and2_1 _21699_ (.A(_03278_),
    .B(_03424_),
    .X(_03426_));
 sky130_fd_sc_hd__nor2_1 _21700_ (.A(_03425_),
    .B(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__xnor2_2 _21701_ (.A(_03423_),
    .B(_03427_),
    .Y(_03428_));
 sky130_fd_sc_hd__or2_1 _21702_ (.A(_03375_),
    .B(_03410_),
    .X(_03429_));
 sky130_fd_sc_hd__xnor2_2 _21703_ (.A(_03428_),
    .B(_03429_),
    .Y(_03430_));
 sky130_fd_sc_hd__xor2_1 _21704_ (.A(_03420_),
    .B(_03430_),
    .X(_03431_));
 sky130_fd_sc_hd__a2bb2o_1 _21705_ (.A1_N(_03382_),
    .A2_N(_03429_),
    .B1(_03411_),
    .B2(_03403_),
    .X(_03432_));
 sky130_fd_sc_hd__nand2_1 _21706_ (.A(_03431_),
    .B(_03432_),
    .Y(_03433_));
 sky130_fd_sc_hd__or2_1 _21707_ (.A(_03431_),
    .B(_03432_),
    .X(_03434_));
 sky130_fd_sc_hd__and2_1 _21708_ (.A(_03433_),
    .B(_03434_),
    .X(_03435_));
 sky130_fd_sc_hd__nand2_1 _21709_ (.A(_03414_),
    .B(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__or2_1 _21710_ (.A(_03414_),
    .B(_03435_),
    .X(_03437_));
 sky130_fd_sc_hd__and2_2 _21711_ (.A(_03436_),
    .B(_03437_),
    .X(_03438_));
 sky130_fd_sc_hd__or2b_1 _21712_ (.A(_03394_),
    .B_N(_03417_),
    .X(_03439_));
 sky130_fd_sc_hd__a21oi_2 _21713_ (.A1(_03389_),
    .A2(_03392_),
    .B1(_03416_),
    .Y(_03440_));
 sky130_fd_sc_hd__o21ba_1 _21714_ (.A1(_03399_),
    .A2(_03439_),
    .B1_N(_03440_),
    .X(_03441_));
 sky130_fd_sc_hd__xnor2_1 _21715_ (.A(_03438_),
    .B(_03441_),
    .Y(_03442_));
 sky130_fd_sc_hd__mux2_1 _21716_ (.A0(\top_inst.deskew_buff_inst.col_input[82] ),
    .A1(_03442_),
    .S(_06140_),
    .X(_03443_));
 sky130_fd_sc_hd__and2_1 _21717_ (.A(_03311_),
    .B(_03443_),
    .X(_03444_));
 sky130_fd_sc_hd__clkbuf_1 _21718_ (.A(_03444_),
    .X(_00840_));
 sky130_fd_sc_hd__or2b_1 _21719_ (.A(_03441_),
    .B_N(_03438_),
    .X(_03445_));
 sky130_fd_sc_hd__o21bai_1 _21720_ (.A1(_03423_),
    .A2(_03426_),
    .B1_N(_03425_),
    .Y(_03446_));
 sky130_fd_sc_hd__a21oi_2 _21721_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[18] ),
    .A2(_03421_),
    .B1(_03422_),
    .Y(_03447_));
 sky130_fd_sc_hd__xnor2_1 _21722_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[19] ),
    .B(_03376_),
    .Y(_03448_));
 sky130_fd_sc_hd__nor2_1 _21723_ (.A(_03278_),
    .B(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__and2_1 _21724_ (.A(_03278_),
    .B(_03448_),
    .X(_03450_));
 sky130_fd_sc_hd__nor2_1 _21725_ (.A(_03449_),
    .B(_03450_),
    .Y(_03451_));
 sky130_fd_sc_hd__xnor2_2 _21726_ (.A(_03447_),
    .B(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__clkbuf_4 _21727_ (.A(_03375_),
    .X(_03453_));
 sky130_fd_sc_hd__nor2_1 _21728_ (.A(_03453_),
    .B(_03428_),
    .Y(_03454_));
 sky130_fd_sc_hd__xor2_1 _21729_ (.A(_03452_),
    .B(_03454_),
    .X(_03455_));
 sky130_fd_sc_hd__nand2_1 _21730_ (.A(_03446_),
    .B(_03455_),
    .Y(_03456_));
 sky130_fd_sc_hd__or2_1 _21731_ (.A(_03446_),
    .B(_03455_),
    .X(_03457_));
 sky130_fd_sc_hd__nand2_1 _21732_ (.A(_03456_),
    .B(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__a22oi_2 _21733_ (.A1(_03420_),
    .A2(_03430_),
    .B1(_03454_),
    .B2(_03410_),
    .Y(_03459_));
 sky130_fd_sc_hd__nor2_1 _21734_ (.A(_03458_),
    .B(_03459_),
    .Y(_03460_));
 sky130_fd_sc_hd__and2_1 _21735_ (.A(_03458_),
    .B(_03459_),
    .X(_03461_));
 sky130_fd_sc_hd__nor2_2 _21736_ (.A(_03460_),
    .B(_03461_),
    .Y(_03462_));
 sky130_fd_sc_hd__xnor2_2 _21737_ (.A(_03433_),
    .B(_03462_),
    .Y(_03463_));
 sky130_fd_sc_hd__a21oi_1 _21738_ (.A1(_03436_),
    .A2(_03445_),
    .B1(_03463_),
    .Y(_03464_));
 sky130_fd_sc_hd__a31o_1 _21739_ (.A1(_03436_),
    .A2(_03445_),
    .A3(_03463_),
    .B1(_01984_),
    .X(_03465_));
 sky130_fd_sc_hd__o221a_1 _21740_ (.A1(net878),
    .A2(_02491_),
    .B1(_03464_),
    .B2(_03465_),
    .C1(_02962_),
    .X(_00841_));
 sky130_fd_sc_hd__nand2_1 _21741_ (.A(_03438_),
    .B(_03463_),
    .Y(_03466_));
 sky130_fd_sc_hd__nand2_1 _21742_ (.A(_03433_),
    .B(_03436_),
    .Y(_03467_));
 sky130_fd_sc_hd__a32oi_4 _21743_ (.A1(_03438_),
    .A2(_03440_),
    .A3(_03463_),
    .B1(_03467_),
    .B2(_03462_),
    .Y(_03468_));
 sky130_fd_sc_hd__o31ai_4 _21744_ (.A1(_03399_),
    .A2(_03439_),
    .A3(_03466_),
    .B1(_03468_),
    .Y(_03469_));
 sky130_fd_sc_hd__nor2_1 _21745_ (.A(_03375_),
    .B(_03452_),
    .Y(_03470_));
 sky130_fd_sc_hd__nand2_1 _21746_ (.A(_03428_),
    .B(_03470_),
    .Y(_03471_));
 sky130_fd_sc_hd__o21bai_2 _21747_ (.A1(_03447_),
    .A2(_03450_),
    .B1_N(_03449_),
    .Y(_03472_));
 sky130_fd_sc_hd__a21oi_2 _21748_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[19] ),
    .A2(_03421_),
    .B1(_03422_),
    .Y(_03473_));
 sky130_fd_sc_hd__xnor2_1 _21749_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[20] ),
    .B(_03376_),
    .Y(_03474_));
 sky130_fd_sc_hd__nor2_1 _21750_ (.A(_03278_),
    .B(_03474_),
    .Y(_03475_));
 sky130_fd_sc_hd__and2_1 _21751_ (.A(_03278_),
    .B(_03474_),
    .X(_03476_));
 sky130_fd_sc_hd__nor2_1 _21752_ (.A(_03475_),
    .B(_03476_),
    .Y(_03477_));
 sky130_fd_sc_hd__xnor2_2 _21753_ (.A(_03473_),
    .B(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__xor2_1 _21754_ (.A(_03478_),
    .B(_03470_),
    .X(_03479_));
 sky130_fd_sc_hd__xnor2_1 _21755_ (.A(_03472_),
    .B(_03479_),
    .Y(_03480_));
 sky130_fd_sc_hd__a21o_1 _21756_ (.A1(_03456_),
    .A2(_03471_),
    .B1(_03480_),
    .X(_03481_));
 sky130_fd_sc_hd__nand3_1 _21757_ (.A(_03456_),
    .B(_03480_),
    .C(_03471_),
    .Y(_03482_));
 sky130_fd_sc_hd__and2_1 _21758_ (.A(_03481_),
    .B(_03482_),
    .X(_03483_));
 sky130_fd_sc_hd__nand2_1 _21759_ (.A(_03460_),
    .B(_03483_),
    .Y(_03484_));
 sky130_fd_sc_hd__or2_1 _21760_ (.A(_03460_),
    .B(_03483_),
    .X(_03485_));
 sky130_fd_sc_hd__and2_1 _21761_ (.A(_03484_),
    .B(_03485_),
    .X(_03486_));
 sky130_fd_sc_hd__nand2_1 _21762_ (.A(_03469_),
    .B(_03486_),
    .Y(_03487_));
 sky130_fd_sc_hd__or2_1 _21763_ (.A(_03469_),
    .B(_03486_),
    .X(_03488_));
 sky130_fd_sc_hd__a21o_1 _21764_ (.A1(_03487_),
    .A2(_03488_),
    .B1(_05732_),
    .X(_03489_));
 sky130_fd_sc_hd__o211a_1 _21765_ (.A1(net886),
    .A2(_06169_),
    .B1(_03489_),
    .C1(_02909_),
    .X(_00842_));
 sky130_fd_sc_hd__o21bai_1 _21766_ (.A1(_03473_),
    .A2(_03476_),
    .B1_N(_03475_),
    .Y(_03490_));
 sky130_fd_sc_hd__a21oi_2 _21767_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[20] ),
    .A2(_03421_),
    .B1(_03422_),
    .Y(_03491_));
 sky130_fd_sc_hd__xnor2_1 _21768_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[21] ),
    .B(_03122_),
    .Y(_03492_));
 sky130_fd_sc_hd__nor2_1 _21769_ (.A(_03278_),
    .B(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__and2_1 _21770_ (.A(_03246_),
    .B(_03492_),
    .X(_03494_));
 sky130_fd_sc_hd__nor2_1 _21771_ (.A(_03493_),
    .B(_03494_),
    .Y(_03495_));
 sky130_fd_sc_hd__xnor2_2 _21772_ (.A(_03491_),
    .B(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__nor2_1 _21773_ (.A(_03375_),
    .B(_03478_),
    .Y(_03497_));
 sky130_fd_sc_hd__xor2_1 _21774_ (.A(_03496_),
    .B(_03497_),
    .X(_03498_));
 sky130_fd_sc_hd__nand2_1 _21775_ (.A(_03490_),
    .B(_03498_),
    .Y(_03499_));
 sky130_fd_sc_hd__or2_1 _21776_ (.A(_03490_),
    .B(_03498_),
    .X(_03500_));
 sky130_fd_sc_hd__nand2_1 _21777_ (.A(_03499_),
    .B(_03500_),
    .Y(_03501_));
 sky130_fd_sc_hd__a22oi_1 _21778_ (.A1(_03472_),
    .A2(_03479_),
    .B1(_03497_),
    .B2(_03452_),
    .Y(_03502_));
 sky130_fd_sc_hd__nor2_1 _21779_ (.A(_03501_),
    .B(_03502_),
    .Y(_03503_));
 sky130_fd_sc_hd__and2_1 _21780_ (.A(_03501_),
    .B(_03502_),
    .X(_03504_));
 sky130_fd_sc_hd__nor2_1 _21781_ (.A(_03503_),
    .B(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__xnor2_2 _21782_ (.A(_03481_),
    .B(_03505_),
    .Y(_03506_));
 sky130_fd_sc_hd__a21oi_1 _21783_ (.A1(_03484_),
    .A2(_03487_),
    .B1(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__a31o_1 _21784_ (.A1(_03484_),
    .A2(_03487_),
    .A3(_03506_),
    .B1(_01984_),
    .X(_03508_));
 sky130_fd_sc_hd__o221a_1 _21785_ (.A1(net648),
    .A2(_02491_),
    .B1(_03507_),
    .B2(_03508_),
    .C1(_02962_),
    .X(_00843_));
 sky130_fd_sc_hd__a21boi_1 _21786_ (.A1(_03481_),
    .A2(_03484_),
    .B1_N(_03505_),
    .Y(_03509_));
 sky130_fd_sc_hd__a31oi_2 _21787_ (.A1(_03469_),
    .A2(_03486_),
    .A3(_03506_),
    .B1(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__nor2_1 _21788_ (.A(_03375_),
    .B(_03496_),
    .Y(_03511_));
 sky130_fd_sc_hd__nand2_1 _21789_ (.A(_03478_),
    .B(_03511_),
    .Y(_03512_));
 sky130_fd_sc_hd__or2_1 _21790_ (.A(_03279_),
    .B(_03492_),
    .X(_03513_));
 sky130_fd_sc_hd__o21ai_1 _21791_ (.A1(_03491_),
    .A2(_03494_),
    .B1(_03513_),
    .Y(_03514_));
 sky130_fd_sc_hd__a21oi_2 _21792_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[21] ),
    .A2(_03421_),
    .B1(_03422_),
    .Y(_03515_));
 sky130_fd_sc_hd__xnor2_1 _21793_ (.A(_03495_),
    .B(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__xor2_1 _21794_ (.A(_03516_),
    .B(_03511_),
    .X(_03517_));
 sky130_fd_sc_hd__xnor2_1 _21795_ (.A(_03514_),
    .B(_03517_),
    .Y(_03518_));
 sky130_fd_sc_hd__a21o_1 _21796_ (.A1(_03499_),
    .A2(_03512_),
    .B1(_03518_),
    .X(_03519_));
 sky130_fd_sc_hd__nand3_1 _21797_ (.A(_03499_),
    .B(_03518_),
    .C(_03512_),
    .Y(_03520_));
 sky130_fd_sc_hd__and2_1 _21798_ (.A(_03519_),
    .B(_03520_),
    .X(_03521_));
 sky130_fd_sc_hd__or2_1 _21799_ (.A(_03503_),
    .B(_03521_),
    .X(_03522_));
 sky130_fd_sc_hd__nand2_1 _21800_ (.A(_03503_),
    .B(_03521_),
    .Y(_03523_));
 sky130_fd_sc_hd__nand2_1 _21801_ (.A(_03522_),
    .B(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__nor2_1 _21802_ (.A(_05405_),
    .B(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__a22o_1 _21803_ (.A1(\top_inst.deskew_buff_inst.col_input[86] ),
    .A2(_05731_),
    .B1(_03510_),
    .B2(_03525_),
    .X(_03526_));
 sky130_fd_sc_hd__and2_1 _21804_ (.A(_03311_),
    .B(_03526_),
    .X(_03527_));
 sky130_fd_sc_hd__clkbuf_1 _21805_ (.A(_03527_),
    .X(_00844_));
 sky130_fd_sc_hd__buf_4 _21806_ (.A(_06168_),
    .X(_03528_));
 sky130_fd_sc_hd__o21ai_1 _21807_ (.A1(_03494_),
    .A2(_03515_),
    .B1(_03513_),
    .Y(_03529_));
 sky130_fd_sc_hd__xnor2_1 _21808_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[23] ),
    .B(_03376_),
    .Y(_03530_));
 sky130_fd_sc_hd__nor2_1 _21809_ (.A(_03278_),
    .B(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__and2_1 _21810_ (.A(_03278_),
    .B(_03530_),
    .X(_03532_));
 sky130_fd_sc_hd__nor2_1 _21811_ (.A(_03531_),
    .B(_03532_),
    .Y(_03533_));
 sky130_fd_sc_hd__xnor2_2 _21812_ (.A(_03515_),
    .B(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__nor2_1 _21813_ (.A(_03375_),
    .B(_03516_),
    .Y(_03535_));
 sky130_fd_sc_hd__xnor2_1 _21814_ (.A(_03534_),
    .B(_03535_),
    .Y(_03536_));
 sky130_fd_sc_hd__xor2_1 _21815_ (.A(_03529_),
    .B(_03536_),
    .X(_03537_));
 sky130_fd_sc_hd__a22oi_1 _21816_ (.A1(_03514_),
    .A2(_03517_),
    .B1(_03535_),
    .B2(_03496_),
    .Y(_03538_));
 sky130_fd_sc_hd__nor2_1 _21817_ (.A(_03537_),
    .B(_03538_),
    .Y(_03539_));
 sky130_fd_sc_hd__and2_1 _21818_ (.A(_03537_),
    .B(_03538_),
    .X(_03540_));
 sky130_fd_sc_hd__nor2_1 _21819_ (.A(_03539_),
    .B(_03540_),
    .Y(_03541_));
 sky130_fd_sc_hd__xnor2_2 _21820_ (.A(_03519_),
    .B(_03541_),
    .Y(_03542_));
 sky130_fd_sc_hd__a21oi_1 _21821_ (.A1(_03510_),
    .A2(_03523_),
    .B1(_03542_),
    .Y(_03543_));
 sky130_fd_sc_hd__a31o_1 _21822_ (.A1(_03510_),
    .A2(_03523_),
    .A3(_03542_),
    .B1(_01984_),
    .X(_03544_));
 sky130_fd_sc_hd__o221a_1 _21823_ (.A1(net670),
    .A2(_03528_),
    .B1(_03543_),
    .B2(_03544_),
    .C1(_02962_),
    .X(_00845_));
 sky130_fd_sc_hd__inv_2 _21824_ (.A(_03524_),
    .Y(_03545_));
 sky130_fd_sc_hd__and4_1 _21825_ (.A(_03486_),
    .B(_03506_),
    .C(_03545_),
    .D(_03542_),
    .X(_03546_));
 sky130_fd_sc_hd__nand2_1 _21826_ (.A(_03519_),
    .B(_03523_),
    .Y(_03547_));
 sky130_fd_sc_hd__a32o_1 _21827_ (.A1(_03509_),
    .A2(_03545_),
    .A3(_03542_),
    .B1(_03547_),
    .B2(_03541_),
    .X(_03548_));
 sky130_fd_sc_hd__a21o_1 _21828_ (.A1(_03469_),
    .A2(_03546_),
    .B1(_03548_),
    .X(_03549_));
 sky130_fd_sc_hd__and2b_1 _21829_ (.A_N(_03536_),
    .B(_03529_),
    .X(_03550_));
 sky130_fd_sc_hd__nor2_1 _21830_ (.A(_03375_),
    .B(_03534_),
    .Y(_03551_));
 sky130_fd_sc_hd__and2_1 _21831_ (.A(_03516_),
    .B(_03551_),
    .X(_03552_));
 sky130_fd_sc_hd__a21o_1 _21832_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[21] ),
    .A2(_03421_),
    .B1(_03422_),
    .X(_03553_));
 sky130_fd_sc_hd__a21o_1 _21833_ (.A1(_03553_),
    .A2(_03533_),
    .B1(_03531_),
    .X(_03554_));
 sky130_fd_sc_hd__a21oi_2 _21834_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[23] ),
    .A2(_03421_),
    .B1(_03422_),
    .Y(_03555_));
 sky130_fd_sc_hd__xnor2_1 _21835_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[24] ),
    .B(_03376_),
    .Y(_03556_));
 sky130_fd_sc_hd__nor2_1 _21836_ (.A(_03279_),
    .B(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__and2_1 _21837_ (.A(_03279_),
    .B(_03556_),
    .X(_03558_));
 sky130_fd_sc_hd__nor2_1 _21838_ (.A(_03557_),
    .B(_03558_),
    .Y(_03559_));
 sky130_fd_sc_hd__xnor2_2 _21839_ (.A(_03555_),
    .B(_03559_),
    .Y(_03560_));
 sky130_fd_sc_hd__xnor2_1 _21840_ (.A(_03560_),
    .B(_03551_),
    .Y(_03561_));
 sky130_fd_sc_hd__xnor2_1 _21841_ (.A(_03554_),
    .B(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hd__o21ai_2 _21842_ (.A1(_03550_),
    .A2(_03552_),
    .B1(_03562_),
    .Y(_03563_));
 sky130_fd_sc_hd__or3_1 _21843_ (.A(_03550_),
    .B(_03562_),
    .C(_03552_),
    .X(_03564_));
 sky130_fd_sc_hd__and2_1 _21844_ (.A(_03563_),
    .B(_03564_),
    .X(_03565_));
 sky130_fd_sc_hd__nand2_1 _21845_ (.A(_03539_),
    .B(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__or2_1 _21846_ (.A(_03539_),
    .B(_03565_),
    .X(_03567_));
 sky130_fd_sc_hd__and2_1 _21847_ (.A(_03566_),
    .B(_03567_),
    .X(_03568_));
 sky130_fd_sc_hd__xor2_1 _21848_ (.A(_03549_),
    .B(_03568_),
    .X(_03569_));
 sky130_fd_sc_hd__or2_1 _21849_ (.A(net524),
    .B(_02638_),
    .X(_03570_));
 sky130_fd_sc_hd__o211a_1 _21850_ (.A1(_03070_),
    .A2(_03569_),
    .B1(_03570_),
    .C1(_02909_),
    .X(_00846_));
 sky130_fd_sc_hd__nand2_1 _21851_ (.A(_03549_),
    .B(_03568_),
    .Y(_03571_));
 sky130_fd_sc_hd__o21bai_2 _21852_ (.A1(_03555_),
    .A2(_03558_),
    .B1_N(_03557_),
    .Y(_03572_));
 sky130_fd_sc_hd__xnor2_1 _21853_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[25] ),
    .B(_03376_),
    .Y(_03573_));
 sky130_fd_sc_hd__or2_2 _21854_ (.A(_03246_),
    .B(_03573_),
    .X(_03574_));
 sky130_fd_sc_hd__nand2_1 _21855_ (.A(_03278_),
    .B(_03573_),
    .Y(_03575_));
 sky130_fd_sc_hd__nand2_2 _21856_ (.A(_03574_),
    .B(_03575_),
    .Y(_03576_));
 sky130_fd_sc_hd__a21oi_1 _21857_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[24] ),
    .A2(_03421_),
    .B1(_03422_),
    .Y(_03577_));
 sky130_fd_sc_hd__or2_1 _21858_ (.A(_03576_),
    .B(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__nand2_1 _21859_ (.A(_03576_),
    .B(_03577_),
    .Y(_03579_));
 sky130_fd_sc_hd__and2_1 _21860_ (.A(_03578_),
    .B(_03579_),
    .X(_03580_));
 sky130_fd_sc_hd__inv_2 _21861_ (.A(_03580_),
    .Y(_03581_));
 sky130_fd_sc_hd__nor2_1 _21862_ (.A(_03453_),
    .B(_03560_),
    .Y(_03582_));
 sky130_fd_sc_hd__xnor2_1 _21863_ (.A(_03581_),
    .B(_03582_),
    .Y(_03583_));
 sky130_fd_sc_hd__xnor2_1 _21864_ (.A(_03572_),
    .B(_03583_),
    .Y(_03584_));
 sky130_fd_sc_hd__and2b_1 _21865_ (.A_N(_03561_),
    .B(_03554_),
    .X(_03585_));
 sky130_fd_sc_hd__a21oi_1 _21866_ (.A1(_03534_),
    .A2(_03582_),
    .B1(_03585_),
    .Y(_03586_));
 sky130_fd_sc_hd__nor2_1 _21867_ (.A(_03584_),
    .B(_03586_),
    .Y(_03587_));
 sky130_fd_sc_hd__and2_1 _21868_ (.A(_03584_),
    .B(_03586_),
    .X(_03588_));
 sky130_fd_sc_hd__nor2_1 _21869_ (.A(_03587_),
    .B(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__xnor2_1 _21870_ (.A(_03563_),
    .B(_03589_),
    .Y(_03590_));
 sky130_fd_sc_hd__a21oi_1 _21871_ (.A1(_03566_),
    .A2(_03571_),
    .B1(_03590_),
    .Y(_03591_));
 sky130_fd_sc_hd__a31o_1 _21872_ (.A1(_03566_),
    .A2(_03571_),
    .A3(_03590_),
    .B1(_01984_),
    .X(_03592_));
 sky130_fd_sc_hd__o221a_1 _21873_ (.A1(net953),
    .A2(_03528_),
    .B1(_03591_),
    .B2(_03592_),
    .C1(_02962_),
    .X(_00847_));
 sky130_fd_sc_hd__and2_1 _21874_ (.A(_03568_),
    .B(_03590_),
    .X(_03593_));
 sky130_fd_sc_hd__a21boi_1 _21875_ (.A1(_03563_),
    .A2(_03566_),
    .B1_N(_03589_),
    .Y(_03594_));
 sky130_fd_sc_hd__a21oi_1 _21876_ (.A1(_03549_),
    .A2(_03593_),
    .B1(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__a21oi_4 _21877_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[25] ),
    .A2(_03421_),
    .B1(_03422_),
    .Y(_03596_));
 sky130_fd_sc_hd__inv_2 _21878_ (.A(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__xnor2_2 _21879_ (.A(_03576_),
    .B(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hd__nor2_1 _21880_ (.A(_03453_),
    .B(_03580_),
    .Y(_03599_));
 sky130_fd_sc_hd__xnor2_1 _21881_ (.A(_03598_),
    .B(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__a21o_1 _21882_ (.A1(_03574_),
    .A2(_03578_),
    .B1(_03600_),
    .X(_03601_));
 sky130_fd_sc_hd__nand3_1 _21883_ (.A(_03574_),
    .B(_03578_),
    .C(_03600_),
    .Y(_03602_));
 sky130_fd_sc_hd__nand2_1 _21884_ (.A(_03601_),
    .B(_03602_),
    .Y(_03603_));
 sky130_fd_sc_hd__a22o_1 _21885_ (.A1(_03572_),
    .A2(_03583_),
    .B1(_03599_),
    .B2(_03560_),
    .X(_03604_));
 sky130_fd_sc_hd__xnor2_1 _21886_ (.A(_03603_),
    .B(_03604_),
    .Y(_03605_));
 sky130_fd_sc_hd__or2_1 _21887_ (.A(_03587_),
    .B(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__nand2_1 _21888_ (.A(_03587_),
    .B(_03605_),
    .Y(_03607_));
 sky130_fd_sc_hd__and2_1 _21889_ (.A(\top_inst.deskew_buff_inst.col_input[90] ),
    .B(_05325_),
    .X(_03608_));
 sky130_fd_sc_hd__a41o_1 _21890_ (.A1(_05312_),
    .A2(_03595_),
    .A3(_03606_),
    .A4(_03607_),
    .B1(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__and2_1 _21891_ (.A(_03311_),
    .B(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__clkbuf_1 _21892_ (.A(_03610_),
    .X(_00848_));
 sky130_fd_sc_hd__or2b_1 _21893_ (.A(_03603_),
    .B_N(_03604_),
    .X(_03611_));
 sky130_fd_sc_hd__o21a_1 _21894_ (.A1(_03576_),
    .A2(_03596_),
    .B1(_03574_),
    .X(_03612_));
 sky130_fd_sc_hd__xnor2_1 _21895_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[27] ),
    .B(_03376_),
    .Y(_03613_));
 sky130_fd_sc_hd__or2_1 _21896_ (.A(_03279_),
    .B(_03613_),
    .X(_03614_));
 sky130_fd_sc_hd__nand2_1 _21897_ (.A(_03279_),
    .B(_03613_),
    .Y(_03615_));
 sky130_fd_sc_hd__nand2_1 _21898_ (.A(_03614_),
    .B(_03615_),
    .Y(_03616_));
 sky130_fd_sc_hd__xnor2_2 _21899_ (.A(_03596_),
    .B(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__xnor2_1 _21900_ (.A(_03453_),
    .B(_03617_),
    .Y(_03618_));
 sky130_fd_sc_hd__mux2_1 _21901_ (.A0(_03618_),
    .A1(_03617_),
    .S(_03598_),
    .X(_03619_));
 sky130_fd_sc_hd__xnor2_1 _21902_ (.A(_03612_),
    .B(_03619_),
    .Y(_03620_));
 sky130_fd_sc_hd__o31a_1 _21903_ (.A1(_03453_),
    .A2(_03581_),
    .A3(_03598_),
    .B1(_03601_),
    .X(_03621_));
 sky130_fd_sc_hd__nor2_1 _21904_ (.A(_03620_),
    .B(_03621_),
    .Y(_03622_));
 sky130_fd_sc_hd__and2_1 _21905_ (.A(_03620_),
    .B(_03621_),
    .X(_03623_));
 sky130_fd_sc_hd__nor2_1 _21906_ (.A(_03622_),
    .B(_03623_),
    .Y(_03624_));
 sky130_fd_sc_hd__xnor2_1 _21907_ (.A(_03611_),
    .B(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__a21oi_1 _21908_ (.A1(_03595_),
    .A2(_03607_),
    .B1(_03625_),
    .Y(_03626_));
 sky130_fd_sc_hd__a31o_1 _21909_ (.A1(_03595_),
    .A2(_03607_),
    .A3(_03625_),
    .B1(_01984_),
    .X(_03627_));
 sky130_fd_sc_hd__o221a_1 _21910_ (.A1(net682),
    .A2(_03528_),
    .B1(_03626_),
    .B2(_03627_),
    .C1(_02962_),
    .X(_00849_));
 sky130_fd_sc_hd__o21a_1 _21911_ (.A1(_03596_),
    .A2(_03616_),
    .B1(_03614_),
    .X(_03628_));
 sky130_fd_sc_hd__or2b_1 _21912_ (.A(_03453_),
    .B_N(_03617_),
    .X(_03629_));
 sky130_fd_sc_hd__a21oi_1 _21913_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[27] ),
    .A2(_03421_),
    .B1(_03422_),
    .Y(_03630_));
 sky130_fd_sc_hd__or2_1 _21914_ (.A(_03576_),
    .B(_03630_),
    .X(_03631_));
 sky130_fd_sc_hd__nand2_1 _21915_ (.A(_03576_),
    .B(_03630_),
    .Y(_03632_));
 sky130_fd_sc_hd__and2_1 _21916_ (.A(_03631_),
    .B(_03632_),
    .X(_03633_));
 sky130_fd_sc_hd__xnor2_1 _21917_ (.A(_03629_),
    .B(_03633_),
    .Y(_03634_));
 sky130_fd_sc_hd__or2b_1 _21918_ (.A(_03628_),
    .B_N(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__or2b_1 _21919_ (.A(_03634_),
    .B_N(_03628_),
    .X(_03636_));
 sky130_fd_sc_hd__nand2_1 _21920_ (.A(_03635_),
    .B(_03636_),
    .Y(_03637_));
 sky130_fd_sc_hd__nand2_1 _21921_ (.A(_03598_),
    .B(_03617_),
    .Y(_03638_));
 sky130_fd_sc_hd__o22ai_2 _21922_ (.A1(_03453_),
    .A2(_03638_),
    .B1(_03619_),
    .B2(_03612_),
    .Y(_03639_));
 sky130_fd_sc_hd__xnor2_1 _21923_ (.A(_03637_),
    .B(_03639_),
    .Y(_03640_));
 sky130_fd_sc_hd__nor2_1 _21924_ (.A(_03622_),
    .B(_03640_),
    .Y(_03641_));
 sky130_fd_sc_hd__and3_1 _21925_ (.A(_03606_),
    .B(_03607_),
    .C(_03625_),
    .X(_03642_));
 sky130_fd_sc_hd__and2_1 _21926_ (.A(_03593_),
    .B(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__nand2_1 _21927_ (.A(_03611_),
    .B(_03607_),
    .Y(_03644_));
 sky130_fd_sc_hd__a22o_1 _21928_ (.A1(_03594_),
    .A2(_03642_),
    .B1(_03644_),
    .B2(_03624_),
    .X(_03645_));
 sky130_fd_sc_hd__nand2_1 _21929_ (.A(_03622_),
    .B(_03640_),
    .Y(_03646_));
 sky130_fd_sc_hd__inv_2 _21930_ (.A(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__a211o_1 _21931_ (.A1(_03549_),
    .A2(_03643_),
    .B1(_03645_),
    .C1(_03647_),
    .X(_03648_));
 sky130_fd_sc_hd__o21ai_1 _21932_ (.A1(_03641_),
    .A2(_03648_),
    .B1(_06178_),
    .Y(_03649_));
 sky130_fd_sc_hd__o211a_1 _21933_ (.A1(net668),
    .A2(_06169_),
    .B1(_03649_),
    .C1(_02909_),
    .X(_00850_));
 sky130_fd_sc_hd__or2b_1 _21934_ (.A(_03637_),
    .B_N(_03639_),
    .X(_03650_));
 sky130_fd_sc_hd__mux2_1 _21935_ (.A0(_03618_),
    .A1(_03617_),
    .S(_03633_),
    .X(_03651_));
 sky130_fd_sc_hd__a21o_1 _21936_ (.A1(_03574_),
    .A2(_03631_),
    .B1(_03651_),
    .X(_03652_));
 sky130_fd_sc_hd__nand3_1 _21937_ (.A(_03574_),
    .B(_03631_),
    .C(_03651_),
    .Y(_03653_));
 sky130_fd_sc_hd__and2_1 _21938_ (.A(_03652_),
    .B(_03653_),
    .X(_03654_));
 sky130_fd_sc_hd__o31a_1 _21939_ (.A1(_03453_),
    .A2(_03617_),
    .A3(_03633_),
    .B1(_03635_),
    .X(_03655_));
 sky130_fd_sc_hd__xor2_1 _21940_ (.A(_03654_),
    .B(_03655_),
    .X(_03656_));
 sky130_fd_sc_hd__xnor2_1 _21941_ (.A(_03650_),
    .B(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__xnor2_1 _21942_ (.A(_03648_),
    .B(_03657_),
    .Y(_03658_));
 sky130_fd_sc_hd__or2_1 _21943_ (.A(net561),
    .B(_09804_),
    .X(_03659_));
 sky130_fd_sc_hd__clkbuf_4 _21944_ (.A(_02706_),
    .X(_03660_));
 sky130_fd_sc_hd__o211a_1 _21945_ (.A1(_03070_),
    .A2(_03658_),
    .B1(_03659_),
    .C1(_03660_),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _21946_ (.A0(\top_inst.deskew_buff_inst.col_input[94] ),
    .A1(_03658_),
    .S(_06140_),
    .X(_03661_));
 sky130_fd_sc_hd__and2_1 _21947_ (.A(_03311_),
    .B(_03661_),
    .X(_03662_));
 sky130_fd_sc_hd__clkbuf_1 _21948_ (.A(_03662_),
    .X(_00852_));
 sky130_fd_sc_hd__a21oi_1 _21949_ (.A1(_03549_),
    .A2(_03643_),
    .B1(_03645_),
    .Y(_03663_));
 sky130_fd_sc_hd__a21o_1 _21950_ (.A1(_03650_),
    .A2(_03646_),
    .B1(_03656_),
    .X(_03664_));
 sky130_fd_sc_hd__or2b_1 _21951_ (.A(_03629_),
    .B_N(_03633_),
    .X(_03665_));
 sky130_fd_sc_hd__mux2_1 _21952_ (.A0(_03597_),
    .A1(_03616_),
    .S(_03453_),
    .X(_03666_));
 sky130_fd_sc_hd__xnor2_1 _21953_ (.A(_03628_),
    .B(_03666_),
    .Y(_03667_));
 sky130_fd_sc_hd__xnor2_1 _21954_ (.A(_03630_),
    .B(_03667_),
    .Y(_03668_));
 sky130_fd_sc_hd__a21o_1 _21955_ (.A1(_03665_),
    .A2(_03652_),
    .B1(_03668_),
    .X(_03669_));
 sky130_fd_sc_hd__nand3_1 _21956_ (.A(_03665_),
    .B(_03652_),
    .C(_03668_),
    .Y(_03670_));
 sky130_fd_sc_hd__nand4b_1 _21957_ (.A_N(_03655_),
    .B(_03669_),
    .C(_03670_),
    .D(_03654_),
    .Y(_03671_));
 sky130_fd_sc_hd__nand2_1 _21958_ (.A(_02885_),
    .B(_02883_),
    .Y(_03672_));
 sky130_fd_sc_hd__a21o_1 _21959_ (.A1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[25] ),
    .A2(_03672_),
    .B1(_03078_),
    .X(_03673_));
 sky130_fd_sc_hd__a31o_1 _21960_ (.A1(_03279_),
    .A2(_03453_),
    .A3(_03673_),
    .B1(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[27] ),
    .X(_03674_));
 sky130_fd_sc_hd__xnor2_1 _21961_ (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[31] ),
    .B(_03669_),
    .Y(_03675_));
 sky130_fd_sc_hd__xnor2_1 _21962_ (.A(_03674_),
    .B(_03675_),
    .Y(_03676_));
 sky130_fd_sc_hd__and4_1 _21963_ (.A(_03663_),
    .B(_03664_),
    .C(_03671_),
    .D(_03676_),
    .X(_03677_));
 sky130_fd_sc_hd__a31o_1 _21964_ (.A1(_03663_),
    .A2(_03664_),
    .A3(_03671_),
    .B1(_03676_),
    .X(_03678_));
 sky130_fd_sc_hd__nand2_1 _21965_ (.A(_06178_),
    .B(_03678_),
    .Y(_03679_));
 sky130_fd_sc_hd__o221a_1 _21966_ (.A1(net954),
    .A2(_03528_),
    .B1(_03677_),
    .B2(_03679_),
    .C1(_02962_),
    .X(_00853_));
 sky130_fd_sc_hd__clkbuf_4 _21967_ (.A(\top_inst.grid_inst.data_path_wires[18][0] ),
    .X(_03680_));
 sky130_fd_sc_hd__or2_1 _21968_ (.A(_03680_),
    .B(_02869_),
    .X(_03681_));
 sky130_fd_sc_hd__o211a_1 _21969_ (.A1(_02862_),
    .A2(_02877_),
    .B1(_03681_),
    .C1(_03660_),
    .X(_00854_));
 sky130_fd_sc_hd__clkbuf_4 _21970_ (.A(\top_inst.grid_inst.data_path_wires[18][1] ),
    .X(_03682_));
 sky130_fd_sc_hd__or2_1 _21971_ (.A(_03682_),
    .B(_02869_),
    .X(_03683_));
 sky130_fd_sc_hd__o211a_1 _21972_ (.A1(_02864_),
    .A2(_02877_),
    .B1(_03683_),
    .C1(_03660_),
    .X(_00855_));
 sky130_fd_sc_hd__clkbuf_4 _21973_ (.A(\top_inst.grid_inst.data_path_wires[18][2] ),
    .X(_03684_));
 sky130_fd_sc_hd__or2_1 _21974_ (.A(_03684_),
    .B(_02869_),
    .X(_03685_));
 sky130_fd_sc_hd__o211a_1 _21975_ (.A1(_02866_),
    .A2(_02877_),
    .B1(_03685_),
    .C1(_03660_),
    .X(_00856_));
 sky130_fd_sc_hd__clkbuf_4 _21976_ (.A(\top_inst.grid_inst.data_path_wires[18][3] ),
    .X(_03686_));
 sky130_fd_sc_hd__or2_1 _21977_ (.A(_03686_),
    .B(_02869_),
    .X(_03687_));
 sky130_fd_sc_hd__o211a_1 _21978_ (.A1(_02868_),
    .A2(_02877_),
    .B1(_03687_),
    .C1(_03660_),
    .X(_00857_));
 sky130_fd_sc_hd__buf_2 _21979_ (.A(\top_inst.grid_inst.data_path_wires[18][4] ),
    .X(_03688_));
 sky130_fd_sc_hd__or2_1 _21980_ (.A(_03688_),
    .B(_02869_),
    .X(_03689_));
 sky130_fd_sc_hd__o211a_1 _21981_ (.A1(_02871_),
    .A2(_02877_),
    .B1(_03689_),
    .C1(_03660_),
    .X(_00858_));
 sky130_fd_sc_hd__clkbuf_4 _21982_ (.A(\top_inst.grid_inst.data_path_wires[18][5] ),
    .X(_03690_));
 sky130_fd_sc_hd__buf_4 _21983_ (.A(_06619_),
    .X(_03691_));
 sky130_fd_sc_hd__or2_1 _21984_ (.A(_03690_),
    .B(_03691_),
    .X(_03692_));
 sky130_fd_sc_hd__o211a_1 _21985_ (.A1(_02873_),
    .A2(_02877_),
    .B1(_03692_),
    .C1(_03660_),
    .X(_00859_));
 sky130_fd_sc_hd__clkbuf_4 _21986_ (.A(\top_inst.grid_inst.data_path_wires[18][6] ),
    .X(_03693_));
 sky130_fd_sc_hd__or2_1 _21987_ (.A(_03693_),
    .B(_03691_),
    .X(_03694_));
 sky130_fd_sc_hd__o211a_1 _21988_ (.A1(_02875_),
    .A2(_02877_),
    .B1(_03694_),
    .C1(_03660_),
    .X(_00860_));
 sky130_fd_sc_hd__clkbuf_4 _21989_ (.A(\top_inst.grid_inst.data_path_wires[18][7] ),
    .X(_03695_));
 sky130_fd_sc_hd__or2_1 _21990_ (.A(_03695_),
    .B(_03691_),
    .X(_03696_));
 sky130_fd_sc_hd__o211a_1 _21991_ (.A1(_02878_),
    .A2(_02877_),
    .B1(_03696_),
    .C1(_03660_),
    .X(_00861_));
 sky130_fd_sc_hd__buf_2 _21992_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[0] ),
    .X(_03697_));
 sky130_fd_sc_hd__clkbuf_4 _21993_ (.A(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__or2_1 _21994_ (.A(_03698_),
    .B(_05275_),
    .X(_03699_));
 sky130_fd_sc_hd__o211a_1 _21995_ (.A1(_03680_),
    .A2(_02881_),
    .B1(_03699_),
    .C1(_03660_),
    .X(_00862_));
 sky130_fd_sc_hd__clkbuf_4 _21996_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[1] ),
    .X(_03700_));
 sky130_fd_sc_hd__or2_1 _21997_ (.A(_03700_),
    .B(_05275_),
    .X(_03701_));
 sky130_fd_sc_hd__clkbuf_4 _21998_ (.A(_02706_),
    .X(_03702_));
 sky130_fd_sc_hd__o211a_1 _21999_ (.A1(_03682_),
    .A2(_02881_),
    .B1(_03701_),
    .C1(_03702_),
    .X(_00863_));
 sky130_fd_sc_hd__clkbuf_4 _22000_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[2] ),
    .X(_03703_));
 sky130_fd_sc_hd__or2_1 _22001_ (.A(_03703_),
    .B(_05275_),
    .X(_03704_));
 sky130_fd_sc_hd__o211a_1 _22002_ (.A1(_03684_),
    .A2(_05270_),
    .B1(_03704_),
    .C1(_03702_),
    .X(_00864_));
 sky130_fd_sc_hd__buf_2 _22003_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[3] ),
    .X(_03705_));
 sky130_fd_sc_hd__or2_1 _22004_ (.A(_03705_),
    .B(_05275_),
    .X(_03706_));
 sky130_fd_sc_hd__o211a_1 _22005_ (.A1(_03686_),
    .A2(_05270_),
    .B1(_03706_),
    .C1(_03702_),
    .X(_00865_));
 sky130_fd_sc_hd__buf_2 _22006_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[4] ),
    .X(_03707_));
 sky130_fd_sc_hd__or2_1 _22007_ (.A(_03707_),
    .B(_05275_),
    .X(_03708_));
 sky130_fd_sc_hd__o211a_1 _22008_ (.A1(_03688_),
    .A2(_05270_),
    .B1(_03708_),
    .C1(_03702_),
    .X(_00866_));
 sky130_fd_sc_hd__clkbuf_4 _22009_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[5] ),
    .X(_03709_));
 sky130_fd_sc_hd__or2_1 _22010_ (.A(_03709_),
    .B(_05275_),
    .X(_03710_));
 sky130_fd_sc_hd__o211a_1 _22011_ (.A1(_03690_),
    .A2(_05270_),
    .B1(_03710_),
    .C1(_03702_),
    .X(_00867_));
 sky130_fd_sc_hd__buf_2 _22012_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[6] ),
    .X(_03711_));
 sky130_fd_sc_hd__or2_1 _22013_ (.A(_03711_),
    .B(_05275_),
    .X(_03712_));
 sky130_fd_sc_hd__o211a_1 _22014_ (.A1(_03693_),
    .A2(_05270_),
    .B1(_03712_),
    .C1(_03702_),
    .X(_00868_));
 sky130_fd_sc_hd__clkbuf_4 _22015_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[7] ),
    .X(_03713_));
 sky130_fd_sc_hd__or2_1 _22016_ (.A(_03713_),
    .B(_05275_),
    .X(_03714_));
 sky130_fd_sc_hd__o211a_1 _22017_ (.A1(_03695_),
    .A2(_05270_),
    .B1(_03714_),
    .C1(_03702_),
    .X(_00869_));
 sky130_fd_sc_hd__and3_1 _22018_ (.A(_03698_),
    .B(_03680_),
    .C(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[0] ),
    .X(_03715_));
 sky130_fd_sc_hd__a21oi_1 _22019_ (.A1(_03698_),
    .A2(_03680_),
    .B1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[0] ),
    .Y(_03716_));
 sky130_fd_sc_hd__o21ai_1 _22020_ (.A1(_03715_),
    .A2(_03716_),
    .B1(_06178_),
    .Y(_03717_));
 sky130_fd_sc_hd__o211a_1 _22021_ (.A1(net1014),
    .A2(_06169_),
    .B1(_03717_),
    .C1(_03702_),
    .X(_00870_));
 sky130_fd_sc_hd__a22o_1 _22022_ (.A1(_03682_),
    .A2(_03698_),
    .B1(_03680_),
    .B2(_03700_),
    .X(_03718_));
 sky130_fd_sc_hd__nand4_2 _22023_ (.A(_03700_),
    .B(_03682_),
    .C(_03698_),
    .D(_03680_),
    .Y(_03719_));
 sky130_fd_sc_hd__nand3_1 _22024_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[1] ),
    .B(_03718_),
    .C(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__a21o_1 _22025_ (.A1(_03718_),
    .A2(_03719_),
    .B1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[1] ),
    .X(_03721_));
 sky130_fd_sc_hd__a21o_1 _22026_ (.A1(_03720_),
    .A2(_03721_),
    .B1(_03715_),
    .X(_03722_));
 sky130_fd_sc_hd__nand3_1 _22027_ (.A(_03715_),
    .B(_03720_),
    .C(_03721_),
    .Y(_03723_));
 sky130_fd_sc_hd__a21o_1 _22028_ (.A1(_03722_),
    .A2(_03723_),
    .B1(_05732_),
    .X(_03724_));
 sky130_fd_sc_hd__o211a_1 _22029_ (.A1(net581),
    .A2(_06169_),
    .B1(_03724_),
    .C1(_03702_),
    .X(_00871_));
 sky130_fd_sc_hd__nand2_1 _22030_ (.A(_03703_),
    .B(_03680_),
    .Y(_03725_));
 sky130_fd_sc_hd__a22o_1 _22031_ (.A1(_03700_),
    .A2(_03682_),
    .B1(_03698_),
    .B2(_03684_),
    .X(_03726_));
 sky130_fd_sc_hd__nand4_1 _22032_ (.A(_03684_),
    .B(_03700_),
    .C(_03682_),
    .D(_03698_),
    .Y(_03727_));
 sky130_fd_sc_hd__nand2_1 _22033_ (.A(_03726_),
    .B(_03727_),
    .Y(_03728_));
 sky130_fd_sc_hd__xnor2_1 _22034_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[2] ),
    .B(_03728_),
    .Y(_03729_));
 sky130_fd_sc_hd__nand2_1 _22035_ (.A(_03719_),
    .B(_03720_),
    .Y(_03730_));
 sky130_fd_sc_hd__xnor2_1 _22036_ (.A(_03729_),
    .B(_03730_),
    .Y(_03731_));
 sky130_fd_sc_hd__or2_1 _22037_ (.A(_03725_),
    .B(_03731_),
    .X(_03732_));
 sky130_fd_sc_hd__nand2_1 _22038_ (.A(_03725_),
    .B(_03731_),
    .Y(_03733_));
 sky130_fd_sc_hd__and2_1 _22039_ (.A(_03732_),
    .B(_03733_),
    .X(_03734_));
 sky130_fd_sc_hd__xnor2_1 _22040_ (.A(_03723_),
    .B(_03734_),
    .Y(_03735_));
 sky130_fd_sc_hd__or2_1 _22041_ (.A(net1103),
    .B(_09804_),
    .X(_03736_));
 sky130_fd_sc_hd__o211a_1 _22042_ (.A1(_03070_),
    .A2(_03735_),
    .B1(_03736_),
    .C1(_03702_),
    .X(_00872_));
 sky130_fd_sc_hd__and2b_1 _22043_ (.A_N(_03723_),
    .B(_03734_),
    .X(_03737_));
 sky130_fd_sc_hd__nand2_1 _22044_ (.A(_03729_),
    .B(_03730_),
    .Y(_03738_));
 sky130_fd_sc_hd__a22o_1 _22045_ (.A1(_03703_),
    .A2(_03682_),
    .B1(_03680_),
    .B2(_03705_),
    .X(_03739_));
 sky130_fd_sc_hd__and4_2 _22046_ (.A(_03705_),
    .B(_03703_),
    .C(_03682_),
    .D(_03680_),
    .X(_03740_));
 sky130_fd_sc_hd__inv_2 _22047_ (.A(_03740_),
    .Y(_03741_));
 sky130_fd_sc_hd__nand2_1 _22048_ (.A(_03739_),
    .B(_03741_),
    .Y(_03742_));
 sky130_fd_sc_hd__a22o_1 _22049_ (.A1(_03684_),
    .A2(_03700_),
    .B1(_03698_),
    .B2(_03686_),
    .X(_03743_));
 sky130_fd_sc_hd__nand4_1 _22050_ (.A(_03686_),
    .B(_03684_),
    .C(_03700_),
    .D(_03698_),
    .Y(_03744_));
 sky130_fd_sc_hd__and3_1 _22051_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[3] ),
    .B(_03743_),
    .C(_03744_),
    .X(_03745_));
 sky130_fd_sc_hd__a21oi_1 _22052_ (.A1(_03743_),
    .A2(_03744_),
    .B1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[3] ),
    .Y(_03746_));
 sky130_fd_sc_hd__or2_2 _22053_ (.A(_03745_),
    .B(_03746_),
    .X(_03747_));
 sky130_fd_sc_hd__a21boi_4 _22054_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[2] ),
    .A2(_03726_),
    .B1_N(_03727_),
    .Y(_03748_));
 sky130_fd_sc_hd__xnor2_2 _22055_ (.A(_03747_),
    .B(_03748_),
    .Y(_03749_));
 sky130_fd_sc_hd__xnor2_1 _22056_ (.A(_03742_),
    .B(_03749_),
    .Y(_03750_));
 sky130_fd_sc_hd__a21o_1 _22057_ (.A1(_03738_),
    .A2(_03732_),
    .B1(_03750_),
    .X(_03751_));
 sky130_fd_sc_hd__nand3_1 _22058_ (.A(_03738_),
    .B(_03732_),
    .C(_03750_),
    .Y(_03752_));
 sky130_fd_sc_hd__nand3_1 _22059_ (.A(_03737_),
    .B(_03751_),
    .C(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__a21o_1 _22060_ (.A1(_03751_),
    .A2(_03752_),
    .B1(_03737_),
    .X(_03754_));
 sky130_fd_sc_hd__and2_1 _22061_ (.A(\top_inst.deskew_buff_inst.col_input[99] ),
    .B(_05730_),
    .X(_03755_));
 sky130_fd_sc_hd__a31o_1 _22062_ (.A1(_05312_),
    .A2(_03753_),
    .A3(_03754_),
    .B1(_03755_),
    .X(_03756_));
 sky130_fd_sc_hd__and2_1 _22063_ (.A(_03311_),
    .B(_03756_),
    .X(_03757_));
 sky130_fd_sc_hd__clkbuf_1 _22064_ (.A(_03757_),
    .X(_00873_));
 sky130_fd_sc_hd__a22o_1 _22065_ (.A1(\top_inst.grid_inst.data_path_wires[18][3] ),
    .A2(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[1] ),
    .B1(_03697_),
    .B2(\top_inst.grid_inst.data_path_wires[18][4] ),
    .X(_03758_));
 sky130_fd_sc_hd__nand4_1 _22066_ (.A(_03688_),
    .B(_03686_),
    .C(_03700_),
    .D(_03697_),
    .Y(_03759_));
 sky130_fd_sc_hd__nand2_1 _22067_ (.A(_03758_),
    .B(_03759_),
    .Y(_03760_));
 sky130_fd_sc_hd__xor2_2 _22068_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[4] ),
    .B(_03760_),
    .X(_03761_));
 sky130_fd_sc_hd__xnor2_2 _22069_ (.A(_03740_),
    .B(_03761_),
    .Y(_03762_));
 sky130_fd_sc_hd__a21bo_1 _22070_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[3] ),
    .A2(_03743_),
    .B1_N(_03744_),
    .X(_03763_));
 sky130_fd_sc_hd__xnor2_2 _22071_ (.A(_03762_),
    .B(_03763_),
    .Y(_03764_));
 sky130_fd_sc_hd__nand2_2 _22072_ (.A(_03703_),
    .B(_03684_),
    .Y(_03765_));
 sky130_fd_sc_hd__nand4_1 _22073_ (.A(_03707_),
    .B(_03705_),
    .C(\top_inst.grid_inst.data_path_wires[18][1] ),
    .D(\top_inst.grid_inst.data_path_wires[18][0] ),
    .Y(_03766_));
 sky130_fd_sc_hd__a22o_1 _22074_ (.A1(_03705_),
    .A2(\top_inst.grid_inst.data_path_wires[18][1] ),
    .B1(\top_inst.grid_inst.data_path_wires[18][0] ),
    .B2(_03707_),
    .X(_03767_));
 sky130_fd_sc_hd__nand2_1 _22075_ (.A(_03766_),
    .B(_03767_),
    .Y(_03768_));
 sky130_fd_sc_hd__xor2_2 _22076_ (.A(_03765_),
    .B(_03768_),
    .X(_03769_));
 sky130_fd_sc_hd__xnor2_2 _22077_ (.A(_03764_),
    .B(_03769_),
    .Y(_03770_));
 sky130_fd_sc_hd__inv_2 _22078_ (.A(_03739_),
    .Y(_03771_));
 sky130_fd_sc_hd__o32ai_4 _22079_ (.A1(_03771_),
    .A2(_03740_),
    .A3(_03749_),
    .B1(_03748_),
    .B2(_03747_),
    .Y(_03772_));
 sky130_fd_sc_hd__xnor2_2 _22080_ (.A(_03770_),
    .B(_03772_),
    .Y(_03773_));
 sky130_fd_sc_hd__nand2_1 _22081_ (.A(_03751_),
    .B(_03753_),
    .Y(_03774_));
 sky130_fd_sc_hd__nor2_1 _22082_ (.A(_03773_),
    .B(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__a21o_1 _22083_ (.A1(_03773_),
    .A2(_03774_),
    .B1(_07595_),
    .X(_03776_));
 sky130_fd_sc_hd__o221a_1 _22084_ (.A1(net371),
    .A2(_03528_),
    .B1(_03775_),
    .B2(_03776_),
    .C1(_02962_),
    .X(_00874_));
 sky130_fd_sc_hd__nor2_1 _22085_ (.A(_03753_),
    .B(_03773_),
    .Y(_03777_));
 sky130_fd_sc_hd__and2b_1 _22086_ (.A_N(_03764_),
    .B(_03769_),
    .X(_03778_));
 sky130_fd_sc_hd__nand2_1 _22087_ (.A(_03709_),
    .B(_03680_),
    .Y(_03779_));
 sky130_fd_sc_hd__nand2_1 _22088_ (.A(_03686_),
    .B(_03703_),
    .Y(_03780_));
 sky130_fd_sc_hd__a22o_1 _22089_ (.A1(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[3] ),
    .A2(\top_inst.grid_inst.data_path_wires[18][2] ),
    .B1(\top_inst.grid_inst.data_path_wires[18][1] ),
    .B2(_03707_),
    .X(_03781_));
 sky130_fd_sc_hd__nand4_1 _22090_ (.A(_03707_),
    .B(_03705_),
    .C(_03684_),
    .D(\top_inst.grid_inst.data_path_wires[18][1] ),
    .Y(_03782_));
 sky130_fd_sc_hd__nand2_1 _22091_ (.A(_03781_),
    .B(_03782_),
    .Y(_03783_));
 sky130_fd_sc_hd__xor2_2 _22092_ (.A(_03780_),
    .B(_03783_),
    .X(_03784_));
 sky130_fd_sc_hd__xnor2_2 _22093_ (.A(_03779_),
    .B(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__a21boi_2 _22094_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[4] ),
    .A2(_03758_),
    .B1_N(_03759_),
    .Y(_03786_));
 sky130_fd_sc_hd__o21ai_2 _22095_ (.A1(_03765_),
    .A2(_03768_),
    .B1(_03766_),
    .Y(_03787_));
 sky130_fd_sc_hd__a22o_1 _22096_ (.A1(\top_inst.grid_inst.data_path_wires[18][4] ),
    .A2(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[1] ),
    .B1(_03697_),
    .B2(_03690_),
    .X(_03788_));
 sky130_fd_sc_hd__nand4_1 _22097_ (.A(_03690_),
    .B(_03688_),
    .C(_03700_),
    .D(_03697_),
    .Y(_03789_));
 sky130_fd_sc_hd__nand2_1 _22098_ (.A(_03788_),
    .B(_03789_),
    .Y(_03790_));
 sky130_fd_sc_hd__xor2_2 _22099_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[5] ),
    .B(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__xnor2_2 _22100_ (.A(_03787_),
    .B(_03791_),
    .Y(_03792_));
 sky130_fd_sc_hd__xnor2_2 _22101_ (.A(_03786_),
    .B(_03792_),
    .Y(_03793_));
 sky130_fd_sc_hd__xor2_2 _22102_ (.A(_03785_),
    .B(_03793_),
    .X(_03794_));
 sky130_fd_sc_hd__xor2_2 _22103_ (.A(_03778_),
    .B(_03794_),
    .X(_03795_));
 sky130_fd_sc_hd__nor2_1 _22104_ (.A(_03741_),
    .B(_03761_),
    .Y(_03796_));
 sky130_fd_sc_hd__a21o_1 _22105_ (.A1(_03762_),
    .A2(_03763_),
    .B1(_03796_),
    .X(_03797_));
 sky130_fd_sc_hd__xnor2_2 _22106_ (.A(_03795_),
    .B(_03797_),
    .Y(_03798_));
 sky130_fd_sc_hd__nand2_1 _22107_ (.A(_03770_),
    .B(_03772_),
    .Y(_03799_));
 sky130_fd_sc_hd__o21ai_1 _22108_ (.A1(_03751_),
    .A2(_03773_),
    .B1(_03799_),
    .Y(_03800_));
 sky130_fd_sc_hd__xnor2_1 _22109_ (.A(_03798_),
    .B(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__nand2_1 _22110_ (.A(_03777_),
    .B(_03801_),
    .Y(_03802_));
 sky130_fd_sc_hd__o21a_1 _22111_ (.A1(_03777_),
    .A2(_03801_),
    .B1(_10831_),
    .X(_03803_));
 sky130_fd_sc_hd__a22o_1 _22112_ (.A1(\top_inst.deskew_buff_inst.col_input[101] ),
    .A2(_05731_),
    .B1(_03802_),
    .B2(_03803_),
    .X(_03804_));
 sky130_fd_sc_hd__and2_1 _22113_ (.A(_03311_),
    .B(_03804_),
    .X(_03805_));
 sky130_fd_sc_hd__clkbuf_1 _22114_ (.A(_03805_),
    .X(_00875_));
 sky130_fd_sc_hd__nor2_1 _22115_ (.A(_03799_),
    .B(_03798_),
    .Y(_03806_));
 sky130_fd_sc_hd__nand2_1 _22116_ (.A(_03778_),
    .B(_03794_),
    .Y(_03807_));
 sky130_fd_sc_hd__nand2_1 _22117_ (.A(_03795_),
    .B(_03797_),
    .Y(_03808_));
 sky130_fd_sc_hd__or2b_1 _22118_ (.A(_03791_),
    .B_N(_03787_),
    .X(_03809_));
 sky130_fd_sc_hd__or2b_1 _22119_ (.A(_03786_),
    .B_N(_03792_),
    .X(_03810_));
 sky130_fd_sc_hd__and2_1 _22120_ (.A(_03785_),
    .B(_03793_),
    .X(_03811_));
 sky130_fd_sc_hd__a21boi_1 _22121_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[5] ),
    .A2(_03788_),
    .B1_N(_03789_),
    .Y(_03812_));
 sky130_fd_sc_hd__o21a_1 _22122_ (.A1(_03780_),
    .A2(_03783_),
    .B1(_03782_),
    .X(_03813_));
 sky130_fd_sc_hd__a22o_1 _22123_ (.A1(\top_inst.grid_inst.data_path_wires[18][5] ),
    .A2(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[1] ),
    .B1(_03697_),
    .B2(\top_inst.grid_inst.data_path_wires[18][6] ),
    .X(_03814_));
 sky130_fd_sc_hd__nand4_1 _22124_ (.A(\top_inst.grid_inst.data_path_wires[18][6] ),
    .B(\top_inst.grid_inst.data_path_wires[18][5] ),
    .C(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[1] ),
    .D(_03697_),
    .Y(_03815_));
 sky130_fd_sc_hd__and3_1 _22125_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[6] ),
    .B(_03814_),
    .C(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__a21oi_1 _22126_ (.A1(_03814_),
    .A2(_03815_),
    .B1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[6] ),
    .Y(_03817_));
 sky130_fd_sc_hd__or2_1 _22127_ (.A(_03816_),
    .B(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__xor2_1 _22128_ (.A(_03813_),
    .B(_03818_),
    .X(_03819_));
 sky130_fd_sc_hd__xnor2_1 _22129_ (.A(_03812_),
    .B(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hd__or2b_1 _22130_ (.A(_03779_),
    .B_N(_03784_),
    .X(_03821_));
 sky130_fd_sc_hd__a22oi_1 _22131_ (.A1(_03709_),
    .A2(_03682_),
    .B1(\top_inst.grid_inst.data_path_wires[18][0] ),
    .B2(_03711_),
    .Y(_03822_));
 sky130_fd_sc_hd__and4_1 _22132_ (.A(_03711_),
    .B(_03709_),
    .C(_03682_),
    .D(\top_inst.grid_inst.data_path_wires[18][0] ),
    .X(_03823_));
 sky130_fd_sc_hd__nor2_1 _22133_ (.A(_03822_),
    .B(_03823_),
    .Y(_03824_));
 sky130_fd_sc_hd__a22oi_1 _22134_ (.A1(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[3] ),
    .A2(\top_inst.grid_inst.data_path_wires[18][3] ),
    .B1(\top_inst.grid_inst.data_path_wires[18][2] ),
    .B2(_03707_),
    .Y(_03825_));
 sky130_fd_sc_hd__and4_1 _22135_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[4] ),
    .B(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[3] ),
    .C(\top_inst.grid_inst.data_path_wires[18][3] ),
    .D(\top_inst.grid_inst.data_path_wires[18][2] ),
    .X(_03826_));
 sky130_fd_sc_hd__and4bb_1 _22136_ (.A_N(_03825_),
    .B_N(_03826_),
    .C(_03688_),
    .D(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[2] ),
    .X(_03827_));
 sky130_fd_sc_hd__o2bb2a_1 _22137_ (.A1_N(_03688_),
    .A2_N(_03703_),
    .B1(_03825_),
    .B2(_03826_),
    .X(_03828_));
 sky130_fd_sc_hd__nor2_1 _22138_ (.A(_03827_),
    .B(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__xnor2_1 _22139_ (.A(_03824_),
    .B(_03829_),
    .Y(_03830_));
 sky130_fd_sc_hd__xor2_1 _22140_ (.A(_03821_),
    .B(_03830_),
    .X(_03831_));
 sky130_fd_sc_hd__nand2_1 _22141_ (.A(_03820_),
    .B(_03831_),
    .Y(_03832_));
 sky130_fd_sc_hd__or2_1 _22142_ (.A(_03820_),
    .B(_03831_),
    .X(_03833_));
 sky130_fd_sc_hd__and3_1 _22143_ (.A(_03811_),
    .B(_03832_),
    .C(_03833_),
    .X(_03834_));
 sky130_fd_sc_hd__a21oi_1 _22144_ (.A1(_03832_),
    .A2(_03833_),
    .B1(_03811_),
    .Y(_03835_));
 sky130_fd_sc_hd__a211oi_2 _22145_ (.A1(_03809_),
    .A2(_03810_),
    .B1(_03834_),
    .C1(_03835_),
    .Y(_03836_));
 sky130_fd_sc_hd__o211a_1 _22146_ (.A1(_03834_),
    .A2(_03835_),
    .B1(_03809_),
    .C1(_03810_),
    .X(_03837_));
 sky130_fd_sc_hd__a211o_1 _22147_ (.A1(_03807_),
    .A2(_03808_),
    .B1(_03836_),
    .C1(_03837_),
    .X(_03838_));
 sky130_fd_sc_hd__o211ai_1 _22148_ (.A1(_03836_),
    .A2(_03837_),
    .B1(_03807_),
    .C1(_03808_),
    .Y(_03839_));
 sky130_fd_sc_hd__and3_1 _22149_ (.A(_03806_),
    .B(_03838_),
    .C(_03839_),
    .X(_03840_));
 sky130_fd_sc_hd__a21oi_1 _22150_ (.A1(_03838_),
    .A2(_03839_),
    .B1(_03806_),
    .Y(_03841_));
 sky130_fd_sc_hd__nor2_1 _22151_ (.A(_03840_),
    .B(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__o31a_1 _22152_ (.A1(_03751_),
    .A2(_03773_),
    .A3(_03798_),
    .B1(_03802_),
    .X(_03843_));
 sky130_fd_sc_hd__xnor2_1 _22153_ (.A(_03842_),
    .B(_03843_),
    .Y(_03844_));
 sky130_fd_sc_hd__mux2_1 _22154_ (.A0(\top_inst.deskew_buff_inst.col_input[102] ),
    .A1(_03844_),
    .S(_06140_),
    .X(_03845_));
 sky130_fd_sc_hd__and2_1 _22155_ (.A(_03311_),
    .B(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__clkbuf_1 _22156_ (.A(_03846_),
    .X(_00876_));
 sky130_fd_sc_hd__or2b_1 _22157_ (.A(_03812_),
    .B_N(_03819_),
    .X(_03847_));
 sky130_fd_sc_hd__o21ai_1 _22158_ (.A1(_03813_),
    .A2(_03818_),
    .B1(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__o21ai_1 _22159_ (.A1(_03821_),
    .A2(_03830_),
    .B1(_03832_),
    .Y(_03849_));
 sky130_fd_sc_hd__a21bo_1 _22160_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[6] ),
    .A2(_03814_),
    .B1_N(_03815_),
    .X(_03850_));
 sky130_fd_sc_hd__nor2_1 _22161_ (.A(_03826_),
    .B(_03827_),
    .Y(_03851_));
 sky130_fd_sc_hd__a22o_1 _22162_ (.A1(\top_inst.grid_inst.data_path_wires[18][6] ),
    .A2(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[1] ),
    .B1(_03697_),
    .B2(_03695_),
    .X(_03852_));
 sky130_fd_sc_hd__nand4_1 _22163_ (.A(_03695_),
    .B(_03693_),
    .C(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[1] ),
    .D(_03697_),
    .Y(_03853_));
 sky130_fd_sc_hd__nand2_1 _22164_ (.A(_03852_),
    .B(_03853_),
    .Y(_03854_));
 sky130_fd_sc_hd__xor2_2 _22165_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[7] ),
    .B(_03854_),
    .X(_03855_));
 sky130_fd_sc_hd__xor2_1 _22166_ (.A(_03851_),
    .B(_03855_),
    .X(_03856_));
 sky130_fd_sc_hd__nand2_1 _22167_ (.A(_03850_),
    .B(_03856_),
    .Y(_03857_));
 sky130_fd_sc_hd__or2_1 _22168_ (.A(_03850_),
    .B(_03856_),
    .X(_03858_));
 sky130_fd_sc_hd__nand2_1 _22169_ (.A(_03857_),
    .B(_03858_),
    .Y(_03859_));
 sky130_fd_sc_hd__and2_1 _22170_ (.A(_03824_),
    .B(_03829_),
    .X(_03860_));
 sky130_fd_sc_hd__a22o_1 _22171_ (.A1(\top_inst.grid_inst.data_path_wires[18][4] ),
    .A2(_03705_),
    .B1(_03686_),
    .B2(_03707_),
    .X(_03861_));
 sky130_fd_sc_hd__nand4_1 _22172_ (.A(_03707_),
    .B(_03688_),
    .C(_03705_),
    .D(_03686_),
    .Y(_03862_));
 sky130_fd_sc_hd__nand2_1 _22173_ (.A(_03861_),
    .B(_03862_),
    .Y(_03863_));
 sky130_fd_sc_hd__and2_1 _22174_ (.A(_03690_),
    .B(_03703_),
    .X(_03864_));
 sky130_fd_sc_hd__xor2_1 _22175_ (.A(_03863_),
    .B(_03864_),
    .X(_03865_));
 sky130_fd_sc_hd__nand2_1 _22176_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[5] ),
    .B(_03684_),
    .Y(_03866_));
 sky130_fd_sc_hd__nand2_1 _22177_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[6] ),
    .B(\top_inst.grid_inst.data_path_wires[18][1] ),
    .Y(_03867_));
 sky130_fd_sc_hd__and2b_1 _22178_ (.A_N(\top_inst.grid_inst.data_path_wires[18][0] ),
    .B(_03713_),
    .X(_03868_));
 sky130_fd_sc_hd__xnor2_1 _22179_ (.A(_03867_),
    .B(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__xnor2_1 _22180_ (.A(_03866_),
    .B(_03869_),
    .Y(_03870_));
 sky130_fd_sc_hd__xnor2_1 _22181_ (.A(_03823_),
    .B(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__xor2_1 _22182_ (.A(_03865_),
    .B(_03871_),
    .X(_03872_));
 sky130_fd_sc_hd__xnor2_1 _22183_ (.A(_03860_),
    .B(_03872_),
    .Y(_03873_));
 sky130_fd_sc_hd__xnor2_1 _22184_ (.A(_03859_),
    .B(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__xor2_1 _22185_ (.A(_03849_),
    .B(_03874_),
    .X(_03875_));
 sky130_fd_sc_hd__xnor2_1 _22186_ (.A(_03848_),
    .B(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hd__nor2_1 _22187_ (.A(_03834_),
    .B(_03836_),
    .Y(_03877_));
 sky130_fd_sc_hd__xnor2_1 _22188_ (.A(_03876_),
    .B(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__xnor2_1 _22189_ (.A(_03713_),
    .B(_03878_),
    .Y(_03879_));
 sky130_fd_sc_hd__xor2_1 _22190_ (.A(_03838_),
    .B(_03879_),
    .X(_03880_));
 sky130_fd_sc_hd__o21bai_2 _22191_ (.A1(_03841_),
    .A2(_03843_),
    .B1_N(_03840_),
    .Y(_03881_));
 sky130_fd_sc_hd__nor2_1 _22192_ (.A(_03880_),
    .B(_03881_),
    .Y(_03882_));
 sky130_fd_sc_hd__a21o_1 _22193_ (.A1(_03880_),
    .A2(_03881_),
    .B1(_05353_),
    .X(_03883_));
 sky130_fd_sc_hd__a2bb2o_1 _22194_ (.A1_N(_03882_),
    .A2_N(_03883_),
    .B1(\top_inst.deskew_buff_inst.col_input[103] ),
    .B2(_05354_),
    .X(_03884_));
 sky130_fd_sc_hd__and2_1 _22195_ (.A(_03311_),
    .B(_03884_),
    .X(_03885_));
 sky130_fd_sc_hd__clkbuf_1 _22196_ (.A(_03885_),
    .X(_00877_));
 sky130_fd_sc_hd__nor2_1 _22197_ (.A(_03838_),
    .B(_03879_),
    .Y(_03886_));
 sky130_fd_sc_hd__a21o_2 _22198_ (.A1(_03880_),
    .A2(_03881_),
    .B1(_03886_),
    .X(_03887_));
 sky130_fd_sc_hd__o21ai_2 _22199_ (.A1(_03851_),
    .A2(_03855_),
    .B1(_03857_),
    .Y(_03888_));
 sky130_fd_sc_hd__a21boi_2 _22200_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[7] ),
    .A2(_03852_),
    .B1_N(_03853_),
    .Y(_03889_));
 sky130_fd_sc_hd__a21boi_2 _22201_ (.A1(_03861_),
    .A2(_03864_),
    .B1_N(_03862_),
    .Y(_03890_));
 sky130_fd_sc_hd__and3_1 _22202_ (.A(\top_inst.grid_inst.data_path_wires[18][7] ),
    .B(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[1] ),
    .C(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[0] ),
    .X(_03891_));
 sky130_fd_sc_hd__o21ai_2 _22203_ (.A1(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[1] ),
    .A2(_03697_),
    .B1(\top_inst.grid_inst.data_path_wires[18][7] ),
    .Y(_03892_));
 sky130_fd_sc_hd__nor2_1 _22204_ (.A(_03891_),
    .B(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__buf_4 _22205_ (.A(_03893_),
    .X(_03894_));
 sky130_fd_sc_hd__xnor2_2 _22206_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[8] ),
    .B(_03894_),
    .Y(_03895_));
 sky130_fd_sc_hd__xor2_2 _22207_ (.A(_03890_),
    .B(_03895_),
    .X(_03896_));
 sky130_fd_sc_hd__xnor2_2 _22208_ (.A(_03889_),
    .B(_03896_),
    .Y(_03897_));
 sky130_fd_sc_hd__a22o_1 _22209_ (.A1(_03707_),
    .A2(_03688_),
    .B1(_03705_),
    .B2(_03690_),
    .X(_03898_));
 sky130_fd_sc_hd__nand4_1 _22210_ (.A(_03690_),
    .B(_03707_),
    .C(_03688_),
    .D(_03705_),
    .Y(_03899_));
 sky130_fd_sc_hd__nand2_1 _22211_ (.A(_03898_),
    .B(_03899_),
    .Y(_03900_));
 sky130_fd_sc_hd__and2_1 _22212_ (.A(_03693_),
    .B(_03703_),
    .X(_03901_));
 sky130_fd_sc_hd__xnor2_2 _22213_ (.A(_03900_),
    .B(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__nand2_1 _22214_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[5] ),
    .B(_03686_),
    .Y(_03903_));
 sky130_fd_sc_hd__and2b_1 _22215_ (.A_N(\top_inst.grid_inst.data_path_wires[18][1] ),
    .B(_03713_),
    .X(_03904_));
 sky130_fd_sc_hd__nand2_1 _22216_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[6] ),
    .B(\top_inst.grid_inst.data_path_wires[18][2] ),
    .Y(_03905_));
 sky130_fd_sc_hd__xnor2_2 _22217_ (.A(_03904_),
    .B(_03905_),
    .Y(_03906_));
 sky130_fd_sc_hd__xnor2_2 _22218_ (.A(_03903_),
    .B(_03906_),
    .Y(_03907_));
 sky130_fd_sc_hd__and3_1 _22219_ (.A(_03711_),
    .B(\top_inst.grid_inst.data_path_wires[18][1] ),
    .C(_03868_),
    .X(_03908_));
 sky130_fd_sc_hd__a31o_1 _22220_ (.A1(_03709_),
    .A2(_03684_),
    .A3(_03869_),
    .B1(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__xor2_2 _22221_ (.A(_03907_),
    .B(_03909_),
    .X(_03910_));
 sky130_fd_sc_hd__xor2_2 _22222_ (.A(_03902_),
    .B(_03910_),
    .X(_03911_));
 sky130_fd_sc_hd__nand2_1 _22223_ (.A(_03823_),
    .B(_03870_),
    .Y(_03912_));
 sky130_fd_sc_hd__o21a_1 _22224_ (.A1(_03865_),
    .A2(_03871_),
    .B1(_03912_),
    .X(_03913_));
 sky130_fd_sc_hd__xnor2_2 _22225_ (.A(_03911_),
    .B(_03913_),
    .Y(_03914_));
 sky130_fd_sc_hd__xnor2_2 _22226_ (.A(_03897_),
    .B(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__nand2_1 _22227_ (.A(_03860_),
    .B(_03872_),
    .Y(_03916_));
 sky130_fd_sc_hd__o21a_1 _22228_ (.A1(_03859_),
    .A2(_03873_),
    .B1(_03916_),
    .X(_03917_));
 sky130_fd_sc_hd__xnor2_2 _22229_ (.A(_03915_),
    .B(_03917_),
    .Y(_03918_));
 sky130_fd_sc_hd__xor2_2 _22230_ (.A(_03888_),
    .B(_03918_),
    .X(_03919_));
 sky130_fd_sc_hd__or2b_1 _22231_ (.A(_03874_),
    .B_N(_03849_),
    .X(_03920_));
 sky130_fd_sc_hd__or2b_1 _22232_ (.A(_03875_),
    .B_N(_03848_),
    .X(_03921_));
 sky130_fd_sc_hd__and2_1 _22233_ (.A(_03920_),
    .B(_03921_),
    .X(_03922_));
 sky130_fd_sc_hd__xnor2_2 _22234_ (.A(_03919_),
    .B(_03922_),
    .Y(_03923_));
 sky130_fd_sc_hd__and2b_1 _22235_ (.A_N(_03877_),
    .B(_03876_),
    .X(_03924_));
 sky130_fd_sc_hd__a21oi_2 _22236_ (.A1(_03713_),
    .A2(_03878_),
    .B1(_03924_),
    .Y(_03925_));
 sky130_fd_sc_hd__xor2_2 _22237_ (.A(_03923_),
    .B(_03925_),
    .X(_03926_));
 sky130_fd_sc_hd__xor2_1 _22238_ (.A(_03887_),
    .B(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__or2_1 _22239_ (.A(net817),
    .B(_09804_),
    .X(_03928_));
 sky130_fd_sc_hd__buf_4 _22240_ (.A(_02706_),
    .X(_03929_));
 sky130_fd_sc_hd__o211a_1 _22241_ (.A1(_03070_),
    .A2(_03927_),
    .B1(_03928_),
    .C1(_03929_),
    .X(_00878_));
 sky130_fd_sc_hd__or2_1 _22242_ (.A(_03923_),
    .B(_03925_),
    .X(_03930_));
 sky130_fd_sc_hd__nand2_1 _22243_ (.A(_03887_),
    .B(_03926_),
    .Y(_03931_));
 sky130_fd_sc_hd__or2_2 _22244_ (.A(_03919_),
    .B(_03922_),
    .X(_03932_));
 sky130_fd_sc_hd__or2_1 _22245_ (.A(_03915_),
    .B(_03917_),
    .X(_03933_));
 sky130_fd_sc_hd__or2b_1 _22246_ (.A(_03918_),
    .B_N(_03888_),
    .X(_03934_));
 sky130_fd_sc_hd__or2b_1 _22247_ (.A(_03889_),
    .B_N(_03896_),
    .X(_03935_));
 sky130_fd_sc_hd__o21ai_1 _22248_ (.A1(_03890_),
    .A2(_03895_),
    .B1(_03935_),
    .Y(_03936_));
 sky130_fd_sc_hd__clkbuf_4 _22249_ (.A(_03894_),
    .X(_03937_));
 sky130_fd_sc_hd__clkbuf_4 _22250_ (.A(_03891_),
    .X(_03938_));
 sky130_fd_sc_hd__a21o_1 _22251_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[8] ),
    .A2(_03937_),
    .B1(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__a21bo_1 _22252_ (.A1(_03898_),
    .A2(_03901_),
    .B1_N(_03899_),
    .X(_03940_));
 sky130_fd_sc_hd__nand2_1 _22253_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[9] ),
    .B(_03894_),
    .Y(_03941_));
 sky130_fd_sc_hd__or2_1 _22254_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[9] ),
    .B(_03894_),
    .X(_03942_));
 sky130_fd_sc_hd__nand2_1 _22255_ (.A(_03941_),
    .B(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__xnor2_2 _22256_ (.A(_03940_),
    .B(_03943_),
    .Y(_03944_));
 sky130_fd_sc_hd__xor2_2 _22257_ (.A(_03939_),
    .B(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__a22o_1 _22258_ (.A1(\top_inst.grid_inst.data_path_wires[18][5] ),
    .A2(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[18][6] ),
    .X(_03946_));
 sky130_fd_sc_hd__and4_1 _22259_ (.A(\top_inst.grid_inst.data_path_wires[18][6] ),
    .B(\top_inst.grid_inst.data_path_wires[18][5] ),
    .C(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[4] ),
    .D(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[3] ),
    .X(_03947_));
 sky130_fd_sc_hd__inv_2 _22260_ (.A(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__and2_1 _22261_ (.A(_03946_),
    .B(_03948_),
    .X(_03949_));
 sky130_fd_sc_hd__nand2_4 _22262_ (.A(\top_inst.grid_inst.data_path_wires[18][7] ),
    .B(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[2] ),
    .Y(_03950_));
 sky130_fd_sc_hd__xnor2_2 _22263_ (.A(_03949_),
    .B(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__nand2_1 _22264_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[5] ),
    .B(\top_inst.grid_inst.data_path_wires[18][4] ),
    .Y(_03952_));
 sky130_fd_sc_hd__and2b_1 _22265_ (.A_N(\top_inst.grid_inst.data_path_wires[18][2] ),
    .B(_03713_),
    .X(_03953_));
 sky130_fd_sc_hd__nand2_1 _22266_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[6] ),
    .B(\top_inst.grid_inst.data_path_wires[18][3] ),
    .Y(_03954_));
 sky130_fd_sc_hd__xnor2_2 _22267_ (.A(_03953_),
    .B(_03954_),
    .Y(_03955_));
 sky130_fd_sc_hd__xnor2_2 _22268_ (.A(_03952_),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__and3_1 _22269_ (.A(_03711_),
    .B(\top_inst.grid_inst.data_path_wires[18][2] ),
    .C(_03904_),
    .X(_03957_));
 sky130_fd_sc_hd__a31o_1 _22270_ (.A1(_03709_),
    .A2(_03686_),
    .A3(_03906_),
    .B1(_03957_),
    .X(_03958_));
 sky130_fd_sc_hd__xor2_2 _22271_ (.A(_03956_),
    .B(_03958_),
    .X(_03959_));
 sky130_fd_sc_hd__xnor2_2 _22272_ (.A(_03951_),
    .B(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__and2_1 _22273_ (.A(_03907_),
    .B(_03909_),
    .X(_03961_));
 sky130_fd_sc_hd__a21o_1 _22274_ (.A1(_03902_),
    .A2(_03910_),
    .B1(_03961_),
    .X(_03962_));
 sky130_fd_sc_hd__xnor2_2 _22275_ (.A(_03960_),
    .B(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__xnor2_1 _22276_ (.A(_03945_),
    .B(_03963_),
    .Y(_03964_));
 sky130_fd_sc_hd__and2b_1 _22277_ (.A_N(_03913_),
    .B(_03911_),
    .X(_03965_));
 sky130_fd_sc_hd__a21oi_1 _22278_ (.A1(_03897_),
    .A2(_03914_),
    .B1(_03965_),
    .Y(_03966_));
 sky130_fd_sc_hd__xor2_1 _22279_ (.A(_03964_),
    .B(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__xnor2_1 _22280_ (.A(_03936_),
    .B(_03967_),
    .Y(_03968_));
 sky130_fd_sc_hd__a21oi_2 _22281_ (.A1(_03933_),
    .A2(_03934_),
    .B1(_03968_),
    .Y(_03969_));
 sky130_fd_sc_hd__and3_1 _22282_ (.A(_03933_),
    .B(_03934_),
    .C(_03968_),
    .X(_03970_));
 sky130_fd_sc_hd__nor2_1 _22283_ (.A(_03969_),
    .B(_03970_),
    .Y(_03971_));
 sky130_fd_sc_hd__xnor2_2 _22284_ (.A(_03932_),
    .B(_03971_),
    .Y(_03972_));
 sky130_fd_sc_hd__a21oi_1 _22285_ (.A1(_03930_),
    .A2(_03931_),
    .B1(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__a31o_1 _22286_ (.A1(_03930_),
    .A2(_03931_),
    .A3(_03972_),
    .B1(_06734_),
    .X(_03974_));
 sky130_fd_sc_hd__o221a_1 _22287_ (.A1(net964),
    .A2(_03528_),
    .B1(_03973_),
    .B2(_03974_),
    .C1(_02962_),
    .X(_00879_));
 sky130_fd_sc_hd__nor2_1 _22288_ (.A(_03964_),
    .B(_03966_),
    .Y(_03975_));
 sky130_fd_sc_hd__a21o_1 _22289_ (.A1(_03936_),
    .A2(_03967_),
    .B1(_03975_),
    .X(_03976_));
 sky130_fd_sc_hd__a32o_1 _22290_ (.A1(_03940_),
    .A2(_03941_),
    .A3(_03942_),
    .B1(_03944_),
    .B2(_03939_),
    .X(_03977_));
 sky130_fd_sc_hd__a21o_1 _22291_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[9] ),
    .A2(_03937_),
    .B1(_03938_),
    .X(_03978_));
 sky130_fd_sc_hd__a31o_1 _22292_ (.A1(_03695_),
    .A2(_03703_),
    .A3(_03946_),
    .B1(_03947_),
    .X(_03979_));
 sky130_fd_sc_hd__xnor2_2 _22293_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[10] ),
    .B(_03894_),
    .Y(_03980_));
 sky130_fd_sc_hd__xnor2_2 _22294_ (.A(_03979_),
    .B(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__xnor2_2 _22295_ (.A(_03978_),
    .B(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__and3_1 _22296_ (.A(\top_inst.grid_inst.data_path_wires[18][7] ),
    .B(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[4] ),
    .C(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[3] ),
    .X(_03983_));
 sky130_fd_sc_hd__a22o_1 _22297_ (.A1(\top_inst.grid_inst.data_path_wires[18][6] ),
    .A2(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[4] ),
    .B1(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[3] ),
    .B2(\top_inst.grid_inst.data_path_wires[18][7] ),
    .X(_03984_));
 sky130_fd_sc_hd__a21bo_1 _22298_ (.A1(_03693_),
    .A2(_03983_),
    .B1_N(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__xor2_2 _22299_ (.A(_03950_),
    .B(_03985_),
    .X(_03986_));
 sky130_fd_sc_hd__nand2_1 _22300_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[5] ),
    .B(_03690_),
    .Y(_03987_));
 sky130_fd_sc_hd__and2b_1 _22301_ (.A_N(\top_inst.grid_inst.data_path_wires[18][3] ),
    .B(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[7] ),
    .X(_03988_));
 sky130_fd_sc_hd__nand2_1 _22302_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[6] ),
    .B(\top_inst.grid_inst.data_path_wires[18][4] ),
    .Y(_03989_));
 sky130_fd_sc_hd__xnor2_2 _22303_ (.A(_03988_),
    .B(_03989_),
    .Y(_03990_));
 sky130_fd_sc_hd__xnor2_2 _22304_ (.A(_03987_),
    .B(_03990_),
    .Y(_03991_));
 sky130_fd_sc_hd__and3_1 _22305_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[6] ),
    .B(\top_inst.grid_inst.data_path_wires[18][3] ),
    .C(_03953_),
    .X(_03992_));
 sky130_fd_sc_hd__a31o_1 _22306_ (.A1(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[5] ),
    .A2(_03688_),
    .A3(_03955_),
    .B1(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__xor2_2 _22307_ (.A(_03991_),
    .B(_03993_),
    .X(_03994_));
 sky130_fd_sc_hd__xnor2_2 _22308_ (.A(_03986_),
    .B(_03994_),
    .Y(_03995_));
 sky130_fd_sc_hd__nand2_1 _22309_ (.A(_03956_),
    .B(_03958_),
    .Y(_03996_));
 sky130_fd_sc_hd__a21boi_2 _22310_ (.A1(_03951_),
    .A2(_03959_),
    .B1_N(_03996_),
    .Y(_03997_));
 sky130_fd_sc_hd__xnor2_2 _22311_ (.A(_03995_),
    .B(_03997_),
    .Y(_03998_));
 sky130_fd_sc_hd__xnor2_2 _22312_ (.A(_03982_),
    .B(_03998_),
    .Y(_03999_));
 sky130_fd_sc_hd__and2b_1 _22313_ (.A_N(_03960_),
    .B(_03962_),
    .X(_04000_));
 sky130_fd_sc_hd__a21oi_2 _22314_ (.A1(_03945_),
    .A2(_03963_),
    .B1(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__xor2_2 _22315_ (.A(_03999_),
    .B(_04001_),
    .X(_04002_));
 sky130_fd_sc_hd__xnor2_2 _22316_ (.A(_03977_),
    .B(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__xnor2_2 _22317_ (.A(_03976_),
    .B(_04003_),
    .Y(_04004_));
 sky130_fd_sc_hd__xor2_2 _22318_ (.A(_03969_),
    .B(_04004_),
    .X(_04005_));
 sky130_fd_sc_hd__a21boi_2 _22319_ (.A1(_03932_),
    .A2(_03930_),
    .B1_N(_03971_),
    .Y(_04006_));
 sky130_fd_sc_hd__a31o_1 _22320_ (.A1(_03887_),
    .A2(_03926_),
    .A3(_03972_),
    .B1(_04006_),
    .X(_04007_));
 sky130_fd_sc_hd__nand2_1 _22321_ (.A(_04005_),
    .B(_04007_),
    .Y(_04008_));
 sky130_fd_sc_hd__o21a_1 _22322_ (.A1(_04005_),
    .A2(_04007_),
    .B1(_05311_),
    .X(_04009_));
 sky130_fd_sc_hd__a22o_1 _22323_ (.A1(\top_inst.deskew_buff_inst.col_input[106] ),
    .A2(_05731_),
    .B1(_04008_),
    .B2(_04009_),
    .X(_04010_));
 sky130_fd_sc_hd__and2_1 _22324_ (.A(_03311_),
    .B(_04010_),
    .X(_04011_));
 sky130_fd_sc_hd__clkbuf_1 _22325_ (.A(_04011_),
    .X(_00880_));
 sky130_fd_sc_hd__nand2_1 _22326_ (.A(_03969_),
    .B(_04004_),
    .Y(_04012_));
 sky130_fd_sc_hd__or2b_1 _22327_ (.A(_04003_),
    .B_N(_03976_),
    .X(_04013_));
 sky130_fd_sc_hd__or2b_1 _22328_ (.A(_03980_),
    .B_N(_03979_),
    .X(_04014_));
 sky130_fd_sc_hd__a21bo_1 _22329_ (.A1(_03978_),
    .A2(_03981_),
    .B1_N(_04014_),
    .X(_04015_));
 sky130_fd_sc_hd__a21o_1 _22330_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[10] ),
    .A2(_03894_),
    .B1(_03938_),
    .X(_04016_));
 sky130_fd_sc_hd__a32o_1 _22331_ (.A1(_03695_),
    .A2(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[2] ),
    .A3(_03984_),
    .B1(_03983_),
    .B2(_03693_),
    .X(_04017_));
 sky130_fd_sc_hd__xnor2_1 _22332_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[11] ),
    .B(_03893_),
    .Y(_04018_));
 sky130_fd_sc_hd__xnor2_1 _22333_ (.A(_04017_),
    .B(_04018_),
    .Y(_04019_));
 sky130_fd_sc_hd__and2_1 _22334_ (.A(_04016_),
    .B(_04019_),
    .X(_04020_));
 sky130_fd_sc_hd__nor2_1 _22335_ (.A(_04016_),
    .B(_04019_),
    .Y(_04021_));
 sky130_fd_sc_hd__or2_1 _22336_ (.A(_04020_),
    .B(_04021_),
    .X(_04022_));
 sky130_fd_sc_hd__o21ai_1 _22337_ (.A1(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[4] ),
    .A2(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[3] ),
    .B1(\top_inst.grid_inst.data_path_wires[18][7] ),
    .Y(_04023_));
 sky130_fd_sc_hd__nor2_2 _22338_ (.A(_03983_),
    .B(_04023_),
    .Y(_04024_));
 sky130_fd_sc_hd__xnor2_4 _22339_ (.A(_03950_),
    .B(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__nand2_1 _22340_ (.A(_03693_),
    .B(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[5] ),
    .Y(_04026_));
 sky130_fd_sc_hd__and2b_1 _22341_ (.A_N(\top_inst.grid_inst.data_path_wires[18][4] ),
    .B(_03713_),
    .X(_04027_));
 sky130_fd_sc_hd__nand2_1 _22342_ (.A(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[6] ),
    .B(\top_inst.grid_inst.data_path_wires[18][5] ),
    .Y(_04028_));
 sky130_fd_sc_hd__xnor2_2 _22343_ (.A(_04027_),
    .B(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__xnor2_2 _22344_ (.A(_04026_),
    .B(_04029_),
    .Y(_04030_));
 sky130_fd_sc_hd__and3_1 _22345_ (.A(_03711_),
    .B(\top_inst.grid_inst.data_path_wires[18][4] ),
    .C(_03988_),
    .X(_04031_));
 sky130_fd_sc_hd__a31o_1 _22346_ (.A1(_03709_),
    .A2(_03690_),
    .A3(_03990_),
    .B1(_04031_),
    .X(_04032_));
 sky130_fd_sc_hd__xor2_2 _22347_ (.A(_04030_),
    .B(_04032_),
    .X(_04033_));
 sky130_fd_sc_hd__xnor2_2 _22348_ (.A(_04025_),
    .B(_04033_),
    .Y(_04034_));
 sky130_fd_sc_hd__and2_1 _22349_ (.A(_03991_),
    .B(_03993_),
    .X(_04035_));
 sky130_fd_sc_hd__a21oi_2 _22350_ (.A1(_03986_),
    .A2(_03994_),
    .B1(_04035_),
    .Y(_04036_));
 sky130_fd_sc_hd__xnor2_2 _22351_ (.A(_04034_),
    .B(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__xor2_2 _22352_ (.A(_04022_),
    .B(_04037_),
    .X(_04038_));
 sky130_fd_sc_hd__or2_1 _22353_ (.A(_03995_),
    .B(_03997_),
    .X(_04039_));
 sky130_fd_sc_hd__o21a_1 _22354_ (.A1(_03982_),
    .A2(_03998_),
    .B1(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__xor2_2 _22355_ (.A(_04038_),
    .B(_04040_),
    .X(_04041_));
 sky130_fd_sc_hd__xor2_2 _22356_ (.A(_04015_),
    .B(_04041_),
    .X(_04042_));
 sky130_fd_sc_hd__nor2_1 _22357_ (.A(_03999_),
    .B(_04001_),
    .Y(_04043_));
 sky130_fd_sc_hd__a21oi_2 _22358_ (.A1(_03977_),
    .A2(_04002_),
    .B1(_04043_),
    .Y(_04044_));
 sky130_fd_sc_hd__xor2_2 _22359_ (.A(_04042_),
    .B(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__xnor2_2 _22360_ (.A(_04013_),
    .B(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__a21oi_1 _22361_ (.A1(_04012_),
    .A2(_04008_),
    .B1(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__and3_1 _22362_ (.A(_04012_),
    .B(_04008_),
    .C(_04046_),
    .X(_04048_));
 sky130_fd_sc_hd__or2_1 _22363_ (.A(net711),
    .B(_05316_),
    .X(_04049_));
 sky130_fd_sc_hd__o311a_1 _22364_ (.A1(_09787_),
    .A2(_04047_),
    .A3(_04048_),
    .B1(_04049_),
    .C1(_05352_),
    .X(_00881_));
 sky130_fd_sc_hd__and2_1 _22365_ (.A(_04005_),
    .B(_04046_),
    .X(_04050_));
 sky130_fd_sc_hd__and3_1 _22366_ (.A(_03926_),
    .B(_03972_),
    .C(_04050_),
    .X(_04051_));
 sky130_fd_sc_hd__a21boi_2 _22367_ (.A1(_04013_),
    .A2(_04012_),
    .B1_N(_04045_),
    .Y(_04052_));
 sky130_fd_sc_hd__a221oi_4 _22368_ (.A1(_04006_),
    .A2(_04050_),
    .B1(_04051_),
    .B2(_03887_),
    .C1(_04052_),
    .Y(_04053_));
 sky130_fd_sc_hd__nor2_1 _22369_ (.A(_04042_),
    .B(_04044_),
    .Y(_04054_));
 sky130_fd_sc_hd__or2b_1 _22370_ (.A(_04040_),
    .B_N(_04038_),
    .X(_04055_));
 sky130_fd_sc_hd__or2b_1 _22371_ (.A(_04041_),
    .B_N(_04015_),
    .X(_04056_));
 sky130_fd_sc_hd__or2b_1 _22372_ (.A(_04018_),
    .B_N(_04017_),
    .X(_04057_));
 sky130_fd_sc_hd__a21bo_1 _22373_ (.A1(_04016_),
    .A2(_04019_),
    .B1_N(_04057_),
    .X(_04058_));
 sky130_fd_sc_hd__a21o_1 _22374_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[11] ),
    .A2(_03937_),
    .B1(_03938_),
    .X(_04059_));
 sky130_fd_sc_hd__o21ba_1 _22375_ (.A1(_03950_),
    .A2(_04023_),
    .B1_N(_03983_),
    .X(_04060_));
 sky130_fd_sc_hd__clkbuf_4 _22376_ (.A(_04060_),
    .X(_04061_));
 sky130_fd_sc_hd__xnor2_1 _22377_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[12] ),
    .B(_03894_),
    .Y(_04062_));
 sky130_fd_sc_hd__xor2_1 _22378_ (.A(_04061_),
    .B(_04062_),
    .X(_04063_));
 sky130_fd_sc_hd__and2_1 _22379_ (.A(_04059_),
    .B(_04063_),
    .X(_04064_));
 sky130_fd_sc_hd__nor2_1 _22380_ (.A(_04059_),
    .B(_04063_),
    .Y(_04065_));
 sky130_fd_sc_hd__or2_1 _22381_ (.A(_04064_),
    .B(_04065_),
    .X(_04066_));
 sky130_fd_sc_hd__and2_1 _22382_ (.A(_03695_),
    .B(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[5] ),
    .X(_04067_));
 sky130_fd_sc_hd__and2b_1 _22383_ (.A_N(\top_inst.grid_inst.data_path_wires[18][5] ),
    .B(_03713_),
    .X(_04068_));
 sky130_fd_sc_hd__nand2_1 _22384_ (.A(_03711_),
    .B(\top_inst.grid_inst.data_path_wires[18][6] ),
    .Y(_04069_));
 sky130_fd_sc_hd__xor2_1 _22385_ (.A(_04068_),
    .B(_04069_),
    .X(_04070_));
 sky130_fd_sc_hd__xnor2_1 _22386_ (.A(_04067_),
    .B(_04070_),
    .Y(_04071_));
 sky130_fd_sc_hd__and3_1 _22387_ (.A(_03711_),
    .B(_03690_),
    .C(_04027_),
    .X(_04072_));
 sky130_fd_sc_hd__a31o_1 _22388_ (.A1(_03693_),
    .A2(_03709_),
    .A3(_04029_),
    .B1(_04072_),
    .X(_04073_));
 sky130_fd_sc_hd__xor2_1 _22389_ (.A(_04071_),
    .B(_04073_),
    .X(_04074_));
 sky130_fd_sc_hd__xnor2_1 _22390_ (.A(_04025_),
    .B(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__and2_1 _22391_ (.A(_04030_),
    .B(_04032_),
    .X(_04076_));
 sky130_fd_sc_hd__a21oi_1 _22392_ (.A1(_04025_),
    .A2(_04033_),
    .B1(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hd__xnor2_1 _22393_ (.A(_04075_),
    .B(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hd__xor2_1 _22394_ (.A(_04066_),
    .B(_04078_),
    .X(_04079_));
 sky130_fd_sc_hd__o32a_1 _22395_ (.A1(_04020_),
    .A2(_04021_),
    .A3(_04037_),
    .B1(_04036_),
    .B2(_04034_),
    .X(_04080_));
 sky130_fd_sc_hd__xnor2_1 _22396_ (.A(_04079_),
    .B(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__xnor2_1 _22397_ (.A(_04058_),
    .B(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__a21o_1 _22398_ (.A1(_04055_),
    .A2(_04056_),
    .B1(_04082_),
    .X(_04083_));
 sky130_fd_sc_hd__nand3_1 _22399_ (.A(_04055_),
    .B(_04056_),
    .C(_04082_),
    .Y(_04084_));
 sky130_fd_sc_hd__and2_1 _22400_ (.A(_04083_),
    .B(_04084_),
    .X(_04085_));
 sky130_fd_sc_hd__xor2_1 _22401_ (.A(_04054_),
    .B(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__xnor2_1 _22402_ (.A(_04053_),
    .B(_04086_),
    .Y(_04087_));
 sky130_fd_sc_hd__or2_1 _22403_ (.A(net659),
    .B(_09804_),
    .X(_04088_));
 sky130_fd_sc_hd__o211a_1 _22404_ (.A1(_03070_),
    .A2(_04087_),
    .B1(_04088_),
    .C1(_03929_),
    .X(_00882_));
 sky130_fd_sc_hd__a31o_1 _22405_ (.A1(_04005_),
    .A2(_04007_),
    .A3(_04046_),
    .B1(_04052_),
    .X(_04089_));
 sky130_fd_sc_hd__nand2_1 _22406_ (.A(_04054_),
    .B(_04085_),
    .Y(_04090_));
 sky130_fd_sc_hd__a21bo_1 _22407_ (.A1(_04089_),
    .A2(_04086_),
    .B1_N(_04090_),
    .X(_04091_));
 sky130_fd_sc_hd__clkbuf_4 _22408_ (.A(_04061_),
    .X(_04092_));
 sky130_fd_sc_hd__o21bai_1 _22409_ (.A1(_04092_),
    .A2(_04062_),
    .B1_N(_04064_),
    .Y(_04093_));
 sky130_fd_sc_hd__a21o_1 _22410_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[12] ),
    .A2(_03937_),
    .B1(_03938_),
    .X(_04094_));
 sky130_fd_sc_hd__xnor2_1 _22411_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[13] ),
    .B(_03894_),
    .Y(_04095_));
 sky130_fd_sc_hd__xor2_1 _22412_ (.A(_04060_),
    .B(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__and2_1 _22413_ (.A(_04094_),
    .B(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__nor2_1 _22414_ (.A(_04094_),
    .B(_04096_),
    .Y(_04098_));
 sky130_fd_sc_hd__or2_1 _22415_ (.A(_04097_),
    .B(_04098_),
    .X(_04099_));
 sky130_fd_sc_hd__nand2_2 _22416_ (.A(\top_inst.grid_inst.data_path_wires[18][7] ),
    .B(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[6] ),
    .Y(_04100_));
 sky130_fd_sc_hd__or2b_1 _22417_ (.A(\top_inst.grid_inst.data_path_wires[18][6] ),
    .B_N(_03713_),
    .X(_04101_));
 sky130_fd_sc_hd__xnor2_1 _22418_ (.A(_04100_),
    .B(_04101_),
    .Y(_04102_));
 sky130_fd_sc_hd__xnor2_1 _22419_ (.A(_04067_),
    .B(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__nand2_2 _22420_ (.A(_03695_),
    .B(_03709_),
    .Y(_04104_));
 sky130_fd_sc_hd__and3_1 _22421_ (.A(_03711_),
    .B(_03693_),
    .C(_04068_),
    .X(_04105_));
 sky130_fd_sc_hd__o21bai_1 _22422_ (.A1(_04104_),
    .A2(_04070_),
    .B1_N(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__xor2_1 _22423_ (.A(_04103_),
    .B(_04106_),
    .X(_04107_));
 sky130_fd_sc_hd__xnor2_1 _22424_ (.A(_04025_),
    .B(_04107_),
    .Y(_04108_));
 sky130_fd_sc_hd__and2_1 _22425_ (.A(_04071_),
    .B(_04073_),
    .X(_04109_));
 sky130_fd_sc_hd__a21oi_1 _22426_ (.A1(_04025_),
    .A2(_04074_),
    .B1(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__xnor2_1 _22427_ (.A(_04108_),
    .B(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__xor2_1 _22428_ (.A(_04099_),
    .B(_04111_),
    .X(_04112_));
 sky130_fd_sc_hd__o32a_1 _22429_ (.A1(_04064_),
    .A2(_04065_),
    .A3(_04078_),
    .B1(_04077_),
    .B2(_04075_),
    .X(_04113_));
 sky130_fd_sc_hd__xor2_1 _22430_ (.A(_04112_),
    .B(_04113_),
    .X(_04114_));
 sky130_fd_sc_hd__xor2_1 _22431_ (.A(_04093_),
    .B(_04114_),
    .X(_04115_));
 sky130_fd_sc_hd__and2b_1 _22432_ (.A_N(_04080_),
    .B(_04079_),
    .X(_04116_));
 sky130_fd_sc_hd__a21oi_1 _22433_ (.A1(_04058_),
    .A2(_04081_),
    .B1(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__nor2_1 _22434_ (.A(_04115_),
    .B(_04117_),
    .Y(_04118_));
 sky130_fd_sc_hd__and2_1 _22435_ (.A(_04115_),
    .B(_04117_),
    .X(_04119_));
 sky130_fd_sc_hd__nor2_1 _22436_ (.A(_04118_),
    .B(_04119_),
    .Y(_04120_));
 sky130_fd_sc_hd__xnor2_1 _22437_ (.A(_04083_),
    .B(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__xor2_1 _22438_ (.A(_04091_),
    .B(_04121_),
    .X(_04122_));
 sky130_fd_sc_hd__or2_1 _22439_ (.A(net627),
    .B(_09804_),
    .X(_04123_));
 sky130_fd_sc_hd__o211a_1 _22440_ (.A1(_03070_),
    .A2(_04122_),
    .B1(_04123_),
    .C1(_03929_),
    .X(_00883_));
 sky130_fd_sc_hd__or2b_1 _22441_ (.A(_04113_),
    .B_N(_04112_),
    .X(_04124_));
 sky130_fd_sc_hd__or2b_1 _22442_ (.A(_04114_),
    .B_N(_04093_),
    .X(_04125_));
 sky130_fd_sc_hd__o21bai_1 _22443_ (.A1(_04092_),
    .A2(_04095_),
    .B1_N(_04097_),
    .Y(_04126_));
 sky130_fd_sc_hd__a21o_1 _22444_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[13] ),
    .A2(_03937_),
    .B1(_03938_),
    .X(_04127_));
 sky130_fd_sc_hd__xnor2_1 _22445_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[14] ),
    .B(_03894_),
    .Y(_04128_));
 sky130_fd_sc_hd__nor2_1 _22446_ (.A(_04061_),
    .B(_04128_),
    .Y(_04129_));
 sky130_fd_sc_hd__nand2_1 _22447_ (.A(_04061_),
    .B(_04128_),
    .Y(_04130_));
 sky130_fd_sc_hd__and2b_1 _22448_ (.A_N(_04129_),
    .B(_04130_),
    .X(_04131_));
 sky130_fd_sc_hd__xor2_1 _22449_ (.A(_04127_),
    .B(_04131_),
    .X(_04132_));
 sky130_fd_sc_hd__and2_1 _22450_ (.A(_04103_),
    .B(_04106_),
    .X(_04133_));
 sky130_fd_sc_hd__a21o_1 _22451_ (.A1(_04025_),
    .A2(_04107_),
    .B1(_04133_),
    .X(_04134_));
 sky130_fd_sc_hd__inv_2 _22452_ (.A(_03713_),
    .Y(_04135_));
 sky130_fd_sc_hd__o211ai_4 _22453_ (.A1(_04135_),
    .A2(_03695_),
    .B1(_04104_),
    .C1(_04100_),
    .Y(_04136_));
 sky130_fd_sc_hd__nor2_4 _22454_ (.A(_04025_),
    .B(_04136_),
    .Y(_04137_));
 sky130_fd_sc_hd__or2_1 _22455_ (.A(_04135_),
    .B(_04100_),
    .X(_04138_));
 sky130_fd_sc_hd__o22a_1 _22456_ (.A1(_03693_),
    .A2(_04138_),
    .B1(_04102_),
    .B2(_04104_),
    .X(_04139_));
 sky130_fd_sc_hd__and3_1 _22457_ (.A(_03695_),
    .B(_03711_),
    .C(_03709_),
    .X(_04140_));
 sky130_fd_sc_hd__nor3_1 _22458_ (.A(_04025_),
    .B(_04139_),
    .C(_04140_),
    .Y(_04141_));
 sky130_fd_sc_hd__o211a_1 _22459_ (.A1(_04139_),
    .A2(_04140_),
    .B1(_04025_),
    .C1(_04136_),
    .X(_04142_));
 sky130_fd_sc_hd__or3_1 _22460_ (.A(_04137_),
    .B(_04141_),
    .C(_04142_),
    .X(_04143_));
 sky130_fd_sc_hd__xnor2_1 _22461_ (.A(_04134_),
    .B(_04143_),
    .Y(_04144_));
 sky130_fd_sc_hd__xor2_1 _22462_ (.A(_04132_),
    .B(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__o32a_1 _22463_ (.A1(_04097_),
    .A2(_04098_),
    .A3(_04111_),
    .B1(_04110_),
    .B2(_04108_),
    .X(_04146_));
 sky130_fd_sc_hd__xnor2_1 _22464_ (.A(_04145_),
    .B(_04146_),
    .Y(_04147_));
 sky130_fd_sc_hd__xnor2_1 _22465_ (.A(_04126_),
    .B(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__a21o_1 _22466_ (.A1(_04124_),
    .A2(_04125_),
    .B1(_04148_),
    .X(_04149_));
 sky130_fd_sc_hd__nand3_1 _22467_ (.A(_04124_),
    .B(_04125_),
    .C(_04148_),
    .Y(_04150_));
 sky130_fd_sc_hd__and2_1 _22468_ (.A(_04149_),
    .B(_04150_),
    .X(_04151_));
 sky130_fd_sc_hd__xor2_1 _22469_ (.A(_04118_),
    .B(_04151_),
    .X(_04152_));
 sky130_fd_sc_hd__and2_1 _22470_ (.A(_04086_),
    .B(_04121_),
    .X(_04153_));
 sky130_fd_sc_hd__a21boi_1 _22471_ (.A1(_04083_),
    .A2(_04090_),
    .B1_N(_04120_),
    .Y(_04154_));
 sky130_fd_sc_hd__a21o_1 _22472_ (.A1(_04089_),
    .A2(_04153_),
    .B1(_04154_),
    .X(_04155_));
 sky130_fd_sc_hd__nand2_1 _22473_ (.A(_04152_),
    .B(_04155_),
    .Y(_04156_));
 sky130_fd_sc_hd__o21a_1 _22474_ (.A1(_04152_),
    .A2(_04155_),
    .B1(_05311_),
    .X(_04157_));
 sky130_fd_sc_hd__a22o_1 _22475_ (.A1(\top_inst.deskew_buff_inst.col_input[110] ),
    .A2(_05731_),
    .B1(_04156_),
    .B2(_04157_),
    .X(_04158_));
 sky130_fd_sc_hd__and2_1 _22476_ (.A(_07707_),
    .B(_04158_),
    .X(_04159_));
 sky130_fd_sc_hd__clkbuf_1 _22477_ (.A(_04159_),
    .X(_00884_));
 sky130_fd_sc_hd__nand2_1 _22478_ (.A(_04118_),
    .B(_04151_),
    .Y(_04160_));
 sky130_fd_sc_hd__a21o_1 _22479_ (.A1(_04127_),
    .A2(_04130_),
    .B1(_04129_),
    .X(_04161_));
 sky130_fd_sc_hd__nor2_1 _22480_ (.A(_04137_),
    .B(_04141_),
    .Y(_04162_));
 sky130_fd_sc_hd__buf_4 _22481_ (.A(_03937_),
    .X(_04163_));
 sky130_fd_sc_hd__a21o_1 _22482_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[14] ),
    .A2(_04163_),
    .B1(_03938_),
    .X(_04164_));
 sky130_fd_sc_hd__xnor2_1 _22483_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[15] ),
    .B(_03937_),
    .Y(_04165_));
 sky130_fd_sc_hd__nor2_1 _22484_ (.A(_04061_),
    .B(_04165_),
    .Y(_04166_));
 sky130_fd_sc_hd__nand2_1 _22485_ (.A(_04061_),
    .B(_04165_),
    .Y(_04167_));
 sky130_fd_sc_hd__and2b_1 _22486_ (.A_N(_04166_),
    .B(_04167_),
    .X(_04168_));
 sky130_fd_sc_hd__xor2_1 _22487_ (.A(_04164_),
    .B(_04168_),
    .X(_04169_));
 sky130_fd_sc_hd__xnor2_1 _22488_ (.A(_04162_),
    .B(_04169_),
    .Y(_04170_));
 sky130_fd_sc_hd__and2b_1 _22489_ (.A_N(_04143_),
    .B(_04134_),
    .X(_04171_));
 sky130_fd_sc_hd__a21oi_1 _22490_ (.A1(_04132_),
    .A2(_04144_),
    .B1(_04171_),
    .Y(_04172_));
 sky130_fd_sc_hd__xnor2_1 _22491_ (.A(_04170_),
    .B(_04172_),
    .Y(_04173_));
 sky130_fd_sc_hd__xor2_1 _22492_ (.A(_04161_),
    .B(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__and2b_1 _22493_ (.A_N(_04146_),
    .B(_04145_),
    .X(_04175_));
 sky130_fd_sc_hd__a21oi_1 _22494_ (.A1(_04126_),
    .A2(_04147_),
    .B1(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hd__nor2_1 _22495_ (.A(_04174_),
    .B(_04176_),
    .Y(_04177_));
 sky130_fd_sc_hd__and2_1 _22496_ (.A(_04174_),
    .B(_04176_),
    .X(_04178_));
 sky130_fd_sc_hd__nor2_1 _22497_ (.A(_04177_),
    .B(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__xnor2_1 _22498_ (.A(_04149_),
    .B(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__a21oi_1 _22499_ (.A1(_04160_),
    .A2(_04156_),
    .B1(_04180_),
    .Y(_04181_));
 sky130_fd_sc_hd__and3_1 _22500_ (.A(_04160_),
    .B(_04156_),
    .C(_04180_),
    .X(_04182_));
 sky130_fd_sc_hd__or2_1 _22501_ (.A(net654),
    .B(_05316_),
    .X(_04183_));
 sky130_fd_sc_hd__o311a_1 _22502_ (.A1(_05403_),
    .A2(_04181_),
    .A3(_04182_),
    .B1(_04183_),
    .C1(_05352_),
    .X(_00885_));
 sky130_fd_sc_hd__and2_1 _22503_ (.A(_04152_),
    .B(_04180_),
    .X(_04184_));
 sky130_fd_sc_hd__nand2_1 _22504_ (.A(_04153_),
    .B(_04184_),
    .Y(_04185_));
 sky130_fd_sc_hd__nand2_1 _22505_ (.A(_04154_),
    .B(_04184_),
    .Y(_04186_));
 sky130_fd_sc_hd__a21bo_1 _22506_ (.A1(_04149_),
    .A2(_04160_),
    .B1_N(_04179_),
    .X(_04187_));
 sky130_fd_sc_hd__o211a_1 _22507_ (.A1(_04053_),
    .A2(_04185_),
    .B1(_04186_),
    .C1(_04187_),
    .X(_04188_));
 sky130_fd_sc_hd__nor2_1 _22508_ (.A(_04170_),
    .B(_04172_),
    .Y(_04189_));
 sky130_fd_sc_hd__and2b_1 _22509_ (.A_N(_04173_),
    .B(_04161_),
    .X(_04190_));
 sky130_fd_sc_hd__a21o_1 _22510_ (.A1(_04164_),
    .A2(_04167_),
    .B1(_04166_),
    .X(_04191_));
 sky130_fd_sc_hd__or2_2 _22511_ (.A(_04025_),
    .B(_04136_),
    .X(_04192_));
 sky130_fd_sc_hd__a21o_1 _22512_ (.A1(_04192_),
    .A2(_04169_),
    .B1(_04141_),
    .X(_04193_));
 sky130_fd_sc_hd__a21o_1 _22513_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[15] ),
    .A2(_03937_),
    .B1(_03938_),
    .X(_04194_));
 sky130_fd_sc_hd__xnor2_1 _22514_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[16] ),
    .B(_03894_),
    .Y(_04195_));
 sky130_fd_sc_hd__nor2_1 _22515_ (.A(_04061_),
    .B(_04195_),
    .Y(_04196_));
 sky130_fd_sc_hd__and2_1 _22516_ (.A(_04061_),
    .B(_04195_),
    .X(_04197_));
 sky130_fd_sc_hd__nor2_1 _22517_ (.A(_04196_),
    .B(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__xor2_1 _22518_ (.A(_04194_),
    .B(_04198_),
    .X(_04199_));
 sky130_fd_sc_hd__or2_1 _22519_ (.A(_04137_),
    .B(_04199_),
    .X(_04200_));
 sky130_fd_sc_hd__nand2_1 _22520_ (.A(_04137_),
    .B(_04199_),
    .Y(_04201_));
 sky130_fd_sc_hd__and2_1 _22521_ (.A(_04200_),
    .B(_04201_),
    .X(_04202_));
 sky130_fd_sc_hd__xor2_1 _22522_ (.A(_04193_),
    .B(_04202_),
    .X(_04203_));
 sky130_fd_sc_hd__xnor2_1 _22523_ (.A(_04191_),
    .B(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__o21ai_2 _22524_ (.A1(_04189_),
    .A2(_04190_),
    .B1(_04204_),
    .Y(_04205_));
 sky130_fd_sc_hd__or3_1 _22525_ (.A(_04189_),
    .B(_04190_),
    .C(_04204_),
    .X(_04206_));
 sky130_fd_sc_hd__and2_1 _22526_ (.A(_04205_),
    .B(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__nand2_1 _22527_ (.A(_04177_),
    .B(_04207_),
    .Y(_04208_));
 sky130_fd_sc_hd__or2_1 _22528_ (.A(_04177_),
    .B(_04207_),
    .X(_04209_));
 sky130_fd_sc_hd__and2_1 _22529_ (.A(_04208_),
    .B(_04209_),
    .X(_04210_));
 sky130_fd_sc_hd__or2b_1 _22530_ (.A(_04188_),
    .B_N(_04210_),
    .X(_04211_));
 sky130_fd_sc_hd__or2b_1 _22531_ (.A(_04210_),
    .B_N(_04188_),
    .X(_04212_));
 sky130_fd_sc_hd__a21o_1 _22532_ (.A1(_04211_),
    .A2(_04212_),
    .B1(_05732_),
    .X(_04213_));
 sky130_fd_sc_hd__o211a_1 _22533_ (.A1(net508),
    .A2(_06169_),
    .B1(_04213_),
    .C1(_03929_),
    .X(_00886_));
 sky130_fd_sc_hd__a21o_1 _22534_ (.A1(_04194_),
    .A2(_04198_),
    .B1(_04196_),
    .X(_04214_));
 sky130_fd_sc_hd__clkbuf_4 _22535_ (.A(_04163_),
    .X(_04215_));
 sky130_fd_sc_hd__clkbuf_4 _22536_ (.A(_03938_),
    .X(_04216_));
 sky130_fd_sc_hd__a21o_1 _22537_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[16] ),
    .A2(_04215_),
    .B1(_04216_),
    .X(_04217_));
 sky130_fd_sc_hd__buf_2 _22538_ (.A(_04061_),
    .X(_04218_));
 sky130_fd_sc_hd__xnor2_1 _22539_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[17] ),
    .B(_04163_),
    .Y(_04219_));
 sky130_fd_sc_hd__nor2_1 _22540_ (.A(_04218_),
    .B(_04219_),
    .Y(_04220_));
 sky130_fd_sc_hd__nand2_1 _22541_ (.A(_04218_),
    .B(_04219_),
    .Y(_04221_));
 sky130_fd_sc_hd__and2b_1 _22542_ (.A_N(_04220_),
    .B(_04221_),
    .X(_04222_));
 sky130_fd_sc_hd__xor2_2 _22543_ (.A(_04217_),
    .B(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__xnor2_1 _22544_ (.A(_04200_),
    .B(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__nand2_1 _22545_ (.A(_04214_),
    .B(_04224_),
    .Y(_04225_));
 sky130_fd_sc_hd__or2_1 _22546_ (.A(_04214_),
    .B(_04224_),
    .X(_04226_));
 sky130_fd_sc_hd__nand2_1 _22547_ (.A(_04225_),
    .B(_04226_),
    .Y(_04227_));
 sky130_fd_sc_hd__inv_2 _22548_ (.A(_04202_),
    .Y(_04228_));
 sky130_fd_sc_hd__or2b_1 _22549_ (.A(_04203_),
    .B_N(_04191_),
    .X(_04229_));
 sky130_fd_sc_hd__a21boi_1 _22550_ (.A1(_04193_),
    .A2(_04228_),
    .B1_N(_04229_),
    .Y(_04230_));
 sky130_fd_sc_hd__nor2_1 _22551_ (.A(_04227_),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__and2_1 _22552_ (.A(_04227_),
    .B(_04230_),
    .X(_04232_));
 sky130_fd_sc_hd__or2_1 _22553_ (.A(_04231_),
    .B(_04232_),
    .X(_04233_));
 sky130_fd_sc_hd__xor2_1 _22554_ (.A(_04205_),
    .B(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__a21oi_1 _22555_ (.A1(_04208_),
    .A2(_04211_),
    .B1(_04234_),
    .Y(_04235_));
 sky130_fd_sc_hd__a31o_1 _22556_ (.A1(_04208_),
    .A2(_04211_),
    .A3(_04234_),
    .B1(_06734_),
    .X(_04236_));
 sky130_fd_sc_hd__o221a_1 _22557_ (.A1(net923),
    .A2(_03528_),
    .B1(_04235_),
    .B2(_04236_),
    .C1(_09806_),
    .X(_00887_));
 sky130_fd_sc_hd__nor2_1 _22558_ (.A(_04137_),
    .B(_04223_),
    .Y(_04237_));
 sky130_fd_sc_hd__nand2_1 _22559_ (.A(_04199_),
    .B(_04237_),
    .Y(_04238_));
 sky130_fd_sc_hd__a21o_1 _22560_ (.A1(_04217_),
    .A2(_04221_),
    .B1(_04220_),
    .X(_04239_));
 sky130_fd_sc_hd__a21o_1 _22561_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[17] ),
    .A2(_04215_),
    .B1(_04216_),
    .X(_04240_));
 sky130_fd_sc_hd__xnor2_1 _22562_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[18] ),
    .B(_04163_),
    .Y(_04241_));
 sky130_fd_sc_hd__nor2_1 _22563_ (.A(_04092_),
    .B(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__nand2_1 _22564_ (.A(_04092_),
    .B(_04241_),
    .Y(_04243_));
 sky130_fd_sc_hd__and2b_1 _22565_ (.A_N(_04242_),
    .B(_04243_),
    .X(_04244_));
 sky130_fd_sc_hd__xor2_2 _22566_ (.A(_04240_),
    .B(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__xor2_2 _22567_ (.A(_04245_),
    .B(_04237_),
    .X(_04246_));
 sky130_fd_sc_hd__xnor2_1 _22568_ (.A(_04239_),
    .B(_04246_),
    .Y(_04247_));
 sky130_fd_sc_hd__a21o_1 _22569_ (.A1(_04225_),
    .A2(_04238_),
    .B1(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__nand3_1 _22570_ (.A(_04225_),
    .B(_04247_),
    .C(_04238_),
    .Y(_04249_));
 sky130_fd_sc_hd__and2_1 _22571_ (.A(_04248_),
    .B(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__nand2_1 _22572_ (.A(_04231_),
    .B(_04250_),
    .Y(_04251_));
 sky130_fd_sc_hd__or2_1 _22573_ (.A(_04231_),
    .B(_04250_),
    .X(_04252_));
 sky130_fd_sc_hd__and2_1 _22574_ (.A(_04251_),
    .B(_04252_),
    .X(_04253_));
 sky130_fd_sc_hd__nand2_1 _22575_ (.A(_04210_),
    .B(_04234_),
    .Y(_04254_));
 sky130_fd_sc_hd__a21oi_1 _22576_ (.A1(_04205_),
    .A2(_04208_),
    .B1(_04233_),
    .Y(_04255_));
 sky130_fd_sc_hd__o21ba_1 _22577_ (.A1(_04188_),
    .A2(_04254_),
    .B1_N(_04255_),
    .X(_04256_));
 sky130_fd_sc_hd__xnor2_1 _22578_ (.A(_04253_),
    .B(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__mux2_1 _22579_ (.A0(\top_inst.deskew_buff_inst.col_input[114] ),
    .A1(_04257_),
    .S(_06140_),
    .X(_04258_));
 sky130_fd_sc_hd__and2_1 _22580_ (.A(_07707_),
    .B(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__clkbuf_1 _22581_ (.A(_04259_),
    .X(_00888_));
 sky130_fd_sc_hd__or2b_1 _22582_ (.A(_04256_),
    .B_N(_04253_),
    .X(_04260_));
 sky130_fd_sc_hd__a21o_1 _22583_ (.A1(_04240_),
    .A2(_04243_),
    .B1(_04242_),
    .X(_04261_));
 sky130_fd_sc_hd__a21o_1 _22584_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[18] ),
    .A2(_04215_),
    .B1(_04216_),
    .X(_04262_));
 sky130_fd_sc_hd__xnor2_1 _22585_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[19] ),
    .B(_04163_),
    .Y(_04263_));
 sky130_fd_sc_hd__nor2_1 _22586_ (.A(_04218_),
    .B(_04263_),
    .Y(_04264_));
 sky130_fd_sc_hd__nand2_1 _22587_ (.A(_04092_),
    .B(_04263_),
    .Y(_04265_));
 sky130_fd_sc_hd__and2b_1 _22588_ (.A_N(_04264_),
    .B(_04265_),
    .X(_04266_));
 sky130_fd_sc_hd__xor2_2 _22589_ (.A(_04262_),
    .B(_04266_),
    .X(_04267_));
 sky130_fd_sc_hd__clkbuf_4 _22590_ (.A(_04137_),
    .X(_04268_));
 sky130_fd_sc_hd__nor2_1 _22591_ (.A(_04268_),
    .B(_04245_),
    .Y(_04269_));
 sky130_fd_sc_hd__xor2_1 _22592_ (.A(_04267_),
    .B(_04269_),
    .X(_04270_));
 sky130_fd_sc_hd__nand2_1 _22593_ (.A(_04261_),
    .B(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__or2_1 _22594_ (.A(_04261_),
    .B(_04270_),
    .X(_04272_));
 sky130_fd_sc_hd__nand2_1 _22595_ (.A(_04271_),
    .B(_04272_),
    .Y(_04273_));
 sky130_fd_sc_hd__a22oi_2 _22596_ (.A1(_04239_),
    .A2(_04246_),
    .B1(_04269_),
    .B2(_04223_),
    .Y(_04274_));
 sky130_fd_sc_hd__nor2_1 _22597_ (.A(_04273_),
    .B(_04274_),
    .Y(_04275_));
 sky130_fd_sc_hd__and2_1 _22598_ (.A(_04273_),
    .B(_04274_),
    .X(_04276_));
 sky130_fd_sc_hd__nor2_1 _22599_ (.A(_04275_),
    .B(_04276_),
    .Y(_04277_));
 sky130_fd_sc_hd__xnor2_2 _22600_ (.A(_04248_),
    .B(_04277_),
    .Y(_04278_));
 sky130_fd_sc_hd__a21oi_1 _22601_ (.A1(_04251_),
    .A2(_04260_),
    .B1(_04278_),
    .Y(_04279_));
 sky130_fd_sc_hd__a31o_1 _22602_ (.A1(_04251_),
    .A2(_04260_),
    .A3(_04278_),
    .B1(_06734_),
    .X(_04280_));
 sky130_fd_sc_hd__o221a_1 _22603_ (.A1(net542),
    .A2(_03528_),
    .B1(_04279_),
    .B2(_04280_),
    .C1(_09806_),
    .X(_00889_));
 sky130_fd_sc_hd__nand2_1 _22604_ (.A(_04253_),
    .B(_04278_),
    .Y(_04281_));
 sky130_fd_sc_hd__nand3_1 _22605_ (.A(_04253_),
    .B(_04255_),
    .C(_04278_),
    .Y(_04282_));
 sky130_fd_sc_hd__a21bo_1 _22606_ (.A1(_04248_),
    .A2(_04251_),
    .B1_N(_04277_),
    .X(_04283_));
 sky130_fd_sc_hd__o311ai_4 _22607_ (.A1(_04188_),
    .A2(_04254_),
    .A3(_04281_),
    .B1(_04282_),
    .C1(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__nor2_1 _22608_ (.A(_04268_),
    .B(_04267_),
    .Y(_04285_));
 sky130_fd_sc_hd__nand2_1 _22609_ (.A(_04245_),
    .B(_04285_),
    .Y(_04286_));
 sky130_fd_sc_hd__a21o_1 _22610_ (.A1(_04262_),
    .A2(_04265_),
    .B1(_04264_),
    .X(_04287_));
 sky130_fd_sc_hd__a21o_1 _22611_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[19] ),
    .A2(_04215_),
    .B1(_04216_),
    .X(_04288_));
 sky130_fd_sc_hd__xnor2_1 _22612_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[20] ),
    .B(_04163_),
    .Y(_04289_));
 sky130_fd_sc_hd__nor2_1 _22613_ (.A(_04218_),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__nand2_1 _22614_ (.A(_04218_),
    .B(_04289_),
    .Y(_04291_));
 sky130_fd_sc_hd__and2b_1 _22615_ (.A_N(_04290_),
    .B(_04291_),
    .X(_04292_));
 sky130_fd_sc_hd__xor2_2 _22616_ (.A(_04288_),
    .B(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__xor2_2 _22617_ (.A(_04293_),
    .B(_04285_),
    .X(_04294_));
 sky130_fd_sc_hd__xnor2_1 _22618_ (.A(_04287_),
    .B(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__a21o_1 _22619_ (.A1(_04271_),
    .A2(_04286_),
    .B1(_04295_),
    .X(_04296_));
 sky130_fd_sc_hd__nand3_1 _22620_ (.A(_04271_),
    .B(_04295_),
    .C(_04286_),
    .Y(_04297_));
 sky130_fd_sc_hd__and2_1 _22621_ (.A(_04296_),
    .B(_04297_),
    .X(_04298_));
 sky130_fd_sc_hd__nand2_1 _22622_ (.A(_04275_),
    .B(_04298_),
    .Y(_04299_));
 sky130_fd_sc_hd__or2_1 _22623_ (.A(_04275_),
    .B(_04298_),
    .X(_04300_));
 sky130_fd_sc_hd__and2_1 _22624_ (.A(_04299_),
    .B(_04300_),
    .X(_04301_));
 sky130_fd_sc_hd__nand2_1 _22625_ (.A(_04284_),
    .B(_04301_),
    .Y(_04302_));
 sky130_fd_sc_hd__or2_1 _22626_ (.A(_04284_),
    .B(_04301_),
    .X(_04303_));
 sky130_fd_sc_hd__and2_1 _22627_ (.A(_04302_),
    .B(_04303_),
    .X(_04304_));
 sky130_fd_sc_hd__or2_1 _22628_ (.A(net533),
    .B(_09804_),
    .X(_04305_));
 sky130_fd_sc_hd__o211a_1 _22629_ (.A1(_09787_),
    .A2(_04304_),
    .B1(_04305_),
    .C1(_03929_),
    .X(_00890_));
 sky130_fd_sc_hd__a21o_1 _22630_ (.A1(_04288_),
    .A2(_04291_),
    .B1(_04290_),
    .X(_04306_));
 sky130_fd_sc_hd__a21o_1 _22631_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[20] ),
    .A2(_04163_),
    .B1(_03938_),
    .X(_04307_));
 sky130_fd_sc_hd__xnor2_1 _22632_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[21] ),
    .B(_03937_),
    .Y(_04308_));
 sky130_fd_sc_hd__or2_1 _22633_ (.A(_04061_),
    .B(_04308_),
    .X(_04309_));
 sky130_fd_sc_hd__nand2_1 _22634_ (.A(_04218_),
    .B(_04308_),
    .Y(_04310_));
 sky130_fd_sc_hd__and2_2 _22635_ (.A(_04309_),
    .B(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__xor2_2 _22636_ (.A(_04307_),
    .B(_04311_),
    .X(_04312_));
 sky130_fd_sc_hd__nor2_1 _22637_ (.A(_04137_),
    .B(_04293_),
    .Y(_04313_));
 sky130_fd_sc_hd__xor2_1 _22638_ (.A(_04312_),
    .B(_04313_),
    .X(_04314_));
 sky130_fd_sc_hd__nand2_1 _22639_ (.A(_04306_),
    .B(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hd__or2_1 _22640_ (.A(_04306_),
    .B(_04314_),
    .X(_04316_));
 sky130_fd_sc_hd__nand2_1 _22641_ (.A(_04315_),
    .B(_04316_),
    .Y(_04317_));
 sky130_fd_sc_hd__a22oi_2 _22642_ (.A1(_04287_),
    .A2(_04294_),
    .B1(_04313_),
    .B2(_04267_),
    .Y(_04318_));
 sky130_fd_sc_hd__nor2_1 _22643_ (.A(_04317_),
    .B(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__and2_1 _22644_ (.A(_04317_),
    .B(_04318_),
    .X(_04320_));
 sky130_fd_sc_hd__nor2_1 _22645_ (.A(_04319_),
    .B(_04320_),
    .Y(_04321_));
 sky130_fd_sc_hd__xnor2_2 _22646_ (.A(_04296_),
    .B(_04321_),
    .Y(_04322_));
 sky130_fd_sc_hd__a21oi_1 _22647_ (.A1(_04299_),
    .A2(_04302_),
    .B1(_04322_),
    .Y(_04323_));
 sky130_fd_sc_hd__a31o_1 _22648_ (.A1(_04299_),
    .A2(_04302_),
    .A3(_04322_),
    .B1(_06734_),
    .X(_04324_));
 sky130_fd_sc_hd__o221a_1 _22649_ (.A1(net260),
    .A2(_03528_),
    .B1(_04323_),
    .B2(_04324_),
    .C1(_09806_),
    .X(_00891_));
 sky130_fd_sc_hd__a21boi_1 _22650_ (.A1(_04296_),
    .A2(_04299_),
    .B1_N(_04321_),
    .Y(_04325_));
 sky130_fd_sc_hd__a31oi_2 _22651_ (.A1(_04284_),
    .A2(_04301_),
    .A3(_04322_),
    .B1(_04325_),
    .Y(_04326_));
 sky130_fd_sc_hd__nor2_1 _22652_ (.A(_04137_),
    .B(_04312_),
    .Y(_04327_));
 sky130_fd_sc_hd__nand2_1 _22653_ (.A(_04293_),
    .B(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__a21bo_1 _22654_ (.A1(_04307_),
    .A2(_04310_),
    .B1_N(_04309_),
    .X(_04329_));
 sky130_fd_sc_hd__a21oi_2 _22655_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[21] ),
    .A2(_04215_),
    .B1(_04216_),
    .Y(_04330_));
 sky130_fd_sc_hd__xnor2_2 _22656_ (.A(_04311_),
    .B(_04330_),
    .Y(_04331_));
 sky130_fd_sc_hd__xor2_2 _22657_ (.A(_04331_),
    .B(_04327_),
    .X(_04332_));
 sky130_fd_sc_hd__xnor2_1 _22658_ (.A(_04329_),
    .B(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__a21o_1 _22659_ (.A1(_04315_),
    .A2(_04328_),
    .B1(_04333_),
    .X(_04334_));
 sky130_fd_sc_hd__nand3_1 _22660_ (.A(_04315_),
    .B(_04333_),
    .C(_04328_),
    .Y(_04335_));
 sky130_fd_sc_hd__and2_1 _22661_ (.A(_04334_),
    .B(_04335_),
    .X(_04336_));
 sky130_fd_sc_hd__or2_1 _22662_ (.A(_04319_),
    .B(_04336_),
    .X(_04337_));
 sky130_fd_sc_hd__nand2_1 _22663_ (.A(_04319_),
    .B(_04336_),
    .Y(_04338_));
 sky130_fd_sc_hd__nand2_1 _22664_ (.A(_04337_),
    .B(_04338_),
    .Y(_04339_));
 sky130_fd_sc_hd__nor2_1 _22665_ (.A(_05405_),
    .B(_04339_),
    .Y(_04340_));
 sky130_fd_sc_hd__a22o_1 _22666_ (.A1(\top_inst.deskew_buff_inst.col_input[118] ),
    .A2(_05731_),
    .B1(_04326_),
    .B2(_04340_),
    .X(_04341_));
 sky130_fd_sc_hd__and2_1 _22667_ (.A(_07707_),
    .B(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__clkbuf_1 _22668_ (.A(_04342_),
    .X(_00892_));
 sky130_fd_sc_hd__a21o_1 _22669_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[21] ),
    .A2(_04215_),
    .B1(_04216_),
    .X(_04343_));
 sky130_fd_sc_hd__a21bo_1 _22670_ (.A1(_04310_),
    .A2(_04343_),
    .B1_N(_04309_),
    .X(_04344_));
 sky130_fd_sc_hd__xnor2_1 _22671_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[23] ),
    .B(_04163_),
    .Y(_04345_));
 sky130_fd_sc_hd__nor2_1 _22672_ (.A(_04218_),
    .B(_04345_),
    .Y(_04346_));
 sky130_fd_sc_hd__nand2_1 _22673_ (.A(_04218_),
    .B(_04345_),
    .Y(_04347_));
 sky130_fd_sc_hd__and2b_1 _22674_ (.A_N(_04346_),
    .B(_04347_),
    .X(_04348_));
 sky130_fd_sc_hd__xnor2_2 _22675_ (.A(_04330_),
    .B(_04348_),
    .Y(_04349_));
 sky130_fd_sc_hd__nor2_1 _22676_ (.A(_04137_),
    .B(_04331_),
    .Y(_04350_));
 sky130_fd_sc_hd__xnor2_1 _22677_ (.A(_04349_),
    .B(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__xor2_1 _22678_ (.A(_04344_),
    .B(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__a22oi_2 _22679_ (.A1(_04329_),
    .A2(_04332_),
    .B1(_04350_),
    .B2(_04312_),
    .Y(_04353_));
 sky130_fd_sc_hd__nor2_1 _22680_ (.A(_04352_),
    .B(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__and2_1 _22681_ (.A(_04352_),
    .B(_04353_),
    .X(_04355_));
 sky130_fd_sc_hd__nor2_1 _22682_ (.A(_04354_),
    .B(_04355_),
    .Y(_04356_));
 sky130_fd_sc_hd__xnor2_2 _22683_ (.A(_04334_),
    .B(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__a21oi_1 _22684_ (.A1(_04326_),
    .A2(_04338_),
    .B1(_04357_),
    .Y(_04358_));
 sky130_fd_sc_hd__a31o_1 _22685_ (.A1(_04326_),
    .A2(_04338_),
    .A3(_04357_),
    .B1(_06734_),
    .X(_04359_));
 sky130_fd_sc_hd__o221a_1 _22686_ (.A1(net608),
    .A2(_03528_),
    .B1(_04358_),
    .B2(_04359_),
    .C1(_09806_),
    .X(_00893_));
 sky130_fd_sc_hd__inv_2 _22687_ (.A(_04339_),
    .Y(_04360_));
 sky130_fd_sc_hd__and4_1 _22688_ (.A(_04301_),
    .B(_04322_),
    .C(_04360_),
    .D(_04357_),
    .X(_04361_));
 sky130_fd_sc_hd__nand2_1 _22689_ (.A(_04334_),
    .B(_04338_),
    .Y(_04362_));
 sky130_fd_sc_hd__a32o_1 _22690_ (.A1(_04325_),
    .A2(_04360_),
    .A3(_04357_),
    .B1(_04362_),
    .B2(_04356_),
    .X(_04363_));
 sky130_fd_sc_hd__a21o_1 _22691_ (.A1(_04284_),
    .A2(_04361_),
    .B1(_04363_),
    .X(_04364_));
 sky130_fd_sc_hd__and2b_1 _22692_ (.A_N(_04351_),
    .B(_04344_),
    .X(_04365_));
 sky130_fd_sc_hd__nor2_1 _22693_ (.A(_04268_),
    .B(_04349_),
    .Y(_04366_));
 sky130_fd_sc_hd__and2_1 _22694_ (.A(_04331_),
    .B(_04366_),
    .X(_04367_));
 sky130_fd_sc_hd__a21o_1 _22695_ (.A1(_04343_),
    .A2(_04347_),
    .B1(_04346_),
    .X(_04368_));
 sky130_fd_sc_hd__a21o_1 _22696_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[23] ),
    .A2(_04215_),
    .B1(_04216_),
    .X(_04369_));
 sky130_fd_sc_hd__xnor2_1 _22697_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[24] ),
    .B(_04163_),
    .Y(_04370_));
 sky130_fd_sc_hd__nor2_1 _22698_ (.A(_04092_),
    .B(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__nand2_1 _22699_ (.A(_04092_),
    .B(_04370_),
    .Y(_04372_));
 sky130_fd_sc_hd__and2b_1 _22700_ (.A_N(_04371_),
    .B(_04372_),
    .X(_04373_));
 sky130_fd_sc_hd__xor2_2 _22701_ (.A(_04369_),
    .B(_04373_),
    .X(_04374_));
 sky130_fd_sc_hd__xnor2_1 _22702_ (.A(_04374_),
    .B(_04366_),
    .Y(_04375_));
 sky130_fd_sc_hd__xnor2_1 _22703_ (.A(_04368_),
    .B(_04375_),
    .Y(_04376_));
 sky130_fd_sc_hd__o21ai_2 _22704_ (.A1(_04365_),
    .A2(_04367_),
    .B1(_04376_),
    .Y(_04377_));
 sky130_fd_sc_hd__or3_1 _22705_ (.A(_04365_),
    .B(_04376_),
    .C(_04367_),
    .X(_04378_));
 sky130_fd_sc_hd__and2_1 _22706_ (.A(_04377_),
    .B(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__nand2_1 _22707_ (.A(_04354_),
    .B(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__or2_1 _22708_ (.A(_04354_),
    .B(_04379_),
    .X(_04381_));
 sky130_fd_sc_hd__and2_1 _22709_ (.A(_04380_),
    .B(_04381_),
    .X(_04382_));
 sky130_fd_sc_hd__xor2_1 _22710_ (.A(_04364_),
    .B(_04382_),
    .X(_04383_));
 sky130_fd_sc_hd__or2_1 _22711_ (.A(net441),
    .B(_09804_),
    .X(_04384_));
 sky130_fd_sc_hd__o211a_1 _22712_ (.A1(_09787_),
    .A2(_04383_),
    .B1(_04384_),
    .C1(_03929_),
    .X(_00894_));
 sky130_fd_sc_hd__nand2_1 _22713_ (.A(_04364_),
    .B(_04382_),
    .Y(_04385_));
 sky130_fd_sc_hd__a21o_1 _22714_ (.A1(_04369_),
    .A2(_04372_),
    .B1(_04371_),
    .X(_04386_));
 sky130_fd_sc_hd__xnor2_1 _22715_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[25] ),
    .B(_03937_),
    .Y(_04387_));
 sky130_fd_sc_hd__or2_2 _22716_ (.A(_04218_),
    .B(_04387_),
    .X(_04388_));
 sky130_fd_sc_hd__nand2_1 _22717_ (.A(_04092_),
    .B(_04387_),
    .Y(_04389_));
 sky130_fd_sc_hd__nand2_2 _22718_ (.A(_04388_),
    .B(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__a21oi_1 _22719_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[24] ),
    .A2(_04215_),
    .B1(_04216_),
    .Y(_04391_));
 sky130_fd_sc_hd__or2_1 _22720_ (.A(_04390_),
    .B(_04391_),
    .X(_04392_));
 sky130_fd_sc_hd__nand2_1 _22721_ (.A(_04390_),
    .B(_04391_),
    .Y(_04393_));
 sky130_fd_sc_hd__and2_1 _22722_ (.A(_04392_),
    .B(_04393_),
    .X(_04394_));
 sky130_fd_sc_hd__inv_2 _22723_ (.A(_04394_),
    .Y(_04395_));
 sky130_fd_sc_hd__nor2_1 _22724_ (.A(_04268_),
    .B(_04374_),
    .Y(_04396_));
 sky130_fd_sc_hd__xnor2_1 _22725_ (.A(_04395_),
    .B(_04396_),
    .Y(_04397_));
 sky130_fd_sc_hd__xnor2_1 _22726_ (.A(_04386_),
    .B(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__and2b_1 _22727_ (.A_N(_04375_),
    .B(_04368_),
    .X(_04399_));
 sky130_fd_sc_hd__a21oi_1 _22728_ (.A1(_04349_),
    .A2(_04396_),
    .B1(_04399_),
    .Y(_04400_));
 sky130_fd_sc_hd__nor2_1 _22729_ (.A(_04398_),
    .B(_04400_),
    .Y(_04401_));
 sky130_fd_sc_hd__and2_1 _22730_ (.A(_04398_),
    .B(_04400_),
    .X(_04402_));
 sky130_fd_sc_hd__nor2_1 _22731_ (.A(_04401_),
    .B(_04402_),
    .Y(_04403_));
 sky130_fd_sc_hd__xnor2_1 _22732_ (.A(_04377_),
    .B(_04403_),
    .Y(_04404_));
 sky130_fd_sc_hd__a21oi_1 _22733_ (.A1(_04380_),
    .A2(_04385_),
    .B1(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__a31o_1 _22734_ (.A1(_04380_),
    .A2(_04385_),
    .A3(_04404_),
    .B1(_06734_),
    .X(_04406_));
 sky130_fd_sc_hd__o221a_1 _22735_ (.A1(net777),
    .A2(_05317_),
    .B1(_04405_),
    .B2(_04406_),
    .C1(_09806_),
    .X(_00895_));
 sky130_fd_sc_hd__and2_1 _22736_ (.A(_04382_),
    .B(_04404_),
    .X(_04407_));
 sky130_fd_sc_hd__a21boi_1 _22737_ (.A1(_04377_),
    .A2(_04380_),
    .B1_N(_04403_),
    .Y(_04408_));
 sky130_fd_sc_hd__a21oi_1 _22738_ (.A1(_04364_),
    .A2(_04407_),
    .B1(_04408_),
    .Y(_04409_));
 sky130_fd_sc_hd__a21oi_4 _22739_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[25] ),
    .A2(_04215_),
    .B1(_04216_),
    .Y(_04410_));
 sky130_fd_sc_hd__inv_2 _22740_ (.A(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__xnor2_2 _22741_ (.A(_04390_),
    .B(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__nor2_1 _22742_ (.A(_04268_),
    .B(_04394_),
    .Y(_04413_));
 sky130_fd_sc_hd__xnor2_1 _22743_ (.A(_04412_),
    .B(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__a21o_1 _22744_ (.A1(_04388_),
    .A2(_04392_),
    .B1(_04414_),
    .X(_04415_));
 sky130_fd_sc_hd__nand3_1 _22745_ (.A(_04388_),
    .B(_04392_),
    .C(_04414_),
    .Y(_04416_));
 sky130_fd_sc_hd__nand2_1 _22746_ (.A(_04415_),
    .B(_04416_),
    .Y(_04417_));
 sky130_fd_sc_hd__a22o_1 _22747_ (.A1(_04386_),
    .A2(_04397_),
    .B1(_04413_),
    .B2(_04374_),
    .X(_04418_));
 sky130_fd_sc_hd__xnor2_1 _22748_ (.A(_04417_),
    .B(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__or2_1 _22749_ (.A(_04401_),
    .B(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__nand2_2 _22750_ (.A(_04401_),
    .B(_04419_),
    .Y(_04421_));
 sky130_fd_sc_hd__and2_1 _22751_ (.A(\top_inst.deskew_buff_inst.col_input[122] ),
    .B(_05325_),
    .X(_04422_));
 sky130_fd_sc_hd__a41o_1 _22752_ (.A1(_05312_),
    .A2(_04409_),
    .A3(_04420_),
    .A4(_04421_),
    .B1(_04422_),
    .X(_04423_));
 sky130_fd_sc_hd__and2_1 _22753_ (.A(_07707_),
    .B(_04423_),
    .X(_04424_));
 sky130_fd_sc_hd__clkbuf_1 _22754_ (.A(_04424_),
    .X(_00896_));
 sky130_fd_sc_hd__or2b_1 _22755_ (.A(_04417_),
    .B_N(_04418_),
    .X(_04425_));
 sky130_fd_sc_hd__o21a_1 _22756_ (.A1(_04390_),
    .A2(_04410_),
    .B1(_04388_),
    .X(_04426_));
 sky130_fd_sc_hd__xnor2_1 _22757_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[27] ),
    .B(_04163_),
    .Y(_04427_));
 sky130_fd_sc_hd__or2_1 _22758_ (.A(_04218_),
    .B(_04427_),
    .X(_04428_));
 sky130_fd_sc_hd__nand2_1 _22759_ (.A(_04092_),
    .B(_04427_),
    .Y(_04429_));
 sky130_fd_sc_hd__nand2_2 _22760_ (.A(_04428_),
    .B(_04429_),
    .Y(_04430_));
 sky130_fd_sc_hd__xnor2_4 _22761_ (.A(_04410_),
    .B(_04430_),
    .Y(_04431_));
 sky130_fd_sc_hd__xnor2_1 _22762_ (.A(_04268_),
    .B(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__mux2_1 _22763_ (.A0(_04432_),
    .A1(_04431_),
    .S(_04412_),
    .X(_04433_));
 sky130_fd_sc_hd__nor2_1 _22764_ (.A(_04426_),
    .B(_04433_),
    .Y(_04434_));
 sky130_fd_sc_hd__and2_1 _22765_ (.A(_04426_),
    .B(_04433_),
    .X(_04435_));
 sky130_fd_sc_hd__or2_1 _22766_ (.A(_04434_),
    .B(_04435_),
    .X(_04436_));
 sky130_fd_sc_hd__o31a_1 _22767_ (.A1(_04268_),
    .A2(_04395_),
    .A3(_04412_),
    .B1(_04415_),
    .X(_04437_));
 sky130_fd_sc_hd__nor2_1 _22768_ (.A(_04436_),
    .B(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__and2_1 _22769_ (.A(_04436_),
    .B(_04437_),
    .X(_04439_));
 sky130_fd_sc_hd__nor2_1 _22770_ (.A(_04438_),
    .B(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__xnor2_1 _22771_ (.A(_04425_),
    .B(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__a21oi_1 _22772_ (.A1(_04409_),
    .A2(_04421_),
    .B1(_04441_),
    .Y(_04442_));
 sky130_fd_sc_hd__a31o_1 _22773_ (.A1(_04409_),
    .A2(_04421_),
    .A3(_04441_),
    .B1(_06734_),
    .X(_04443_));
 sky130_fd_sc_hd__o221a_1 _22774_ (.A1(net724),
    .A2(_05317_),
    .B1(_04442_),
    .B2(_04443_),
    .C1(_09806_),
    .X(_00897_));
 sky130_fd_sc_hd__o21a_1 _22775_ (.A1(_04410_),
    .A2(_04430_),
    .B1(_04428_),
    .X(_04444_));
 sky130_fd_sc_hd__a21oi_2 _22776_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[27] ),
    .A2(_04215_),
    .B1(_04216_),
    .Y(_04445_));
 sky130_fd_sc_hd__or2_1 _22777_ (.A(_04390_),
    .B(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__nand2_1 _22778_ (.A(_04390_),
    .B(_04445_),
    .Y(_04447_));
 sky130_fd_sc_hd__and2_1 _22779_ (.A(_04446_),
    .B(_04447_),
    .X(_04448_));
 sky130_fd_sc_hd__nand3_1 _22780_ (.A(_04192_),
    .B(_04431_),
    .C(_04448_),
    .Y(_04449_));
 sky130_fd_sc_hd__a21o_1 _22781_ (.A1(_04192_),
    .A2(_04431_),
    .B1(_04448_),
    .X(_04450_));
 sky130_fd_sc_hd__and2_1 _22782_ (.A(_04449_),
    .B(_04450_),
    .X(_04451_));
 sky130_fd_sc_hd__or2b_1 _22783_ (.A(_04444_),
    .B_N(_04451_),
    .X(_04452_));
 sky130_fd_sc_hd__or2b_1 _22784_ (.A(_04451_),
    .B_N(_04444_),
    .X(_04453_));
 sky130_fd_sc_hd__nand2_1 _22785_ (.A(_04452_),
    .B(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__a31o_1 _22786_ (.A1(_04192_),
    .A2(_04412_),
    .A3(_04431_),
    .B1(_04434_),
    .X(_04455_));
 sky130_fd_sc_hd__xnor2_1 _22787_ (.A(_04454_),
    .B(_04455_),
    .Y(_04456_));
 sky130_fd_sc_hd__nor2_1 _22788_ (.A(_04438_),
    .B(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__and3_1 _22789_ (.A(_04420_),
    .B(_04421_),
    .C(_04441_),
    .X(_04458_));
 sky130_fd_sc_hd__and2_1 _22790_ (.A(_04407_),
    .B(_04458_),
    .X(_04459_));
 sky130_fd_sc_hd__nand2_1 _22791_ (.A(_04425_),
    .B(_04421_),
    .Y(_04460_));
 sky130_fd_sc_hd__a22o_1 _22792_ (.A1(_04408_),
    .A2(_04458_),
    .B1(_04460_),
    .B2(_04440_),
    .X(_04461_));
 sky130_fd_sc_hd__nand2_1 _22793_ (.A(_04438_),
    .B(_04456_),
    .Y(_04462_));
 sky130_fd_sc_hd__inv_2 _22794_ (.A(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__a211o_1 _22795_ (.A1(_04364_),
    .A2(_04459_),
    .B1(_04461_),
    .C1(_04463_),
    .X(_04464_));
 sky130_fd_sc_hd__o21ai_1 _22796_ (.A1(_04457_),
    .A2(_04464_),
    .B1(_06178_),
    .Y(_04465_));
 sky130_fd_sc_hd__o211a_1 _22797_ (.A1(net564),
    .A2(_06169_),
    .B1(_04465_),
    .C1(_03929_),
    .X(_00898_));
 sky130_fd_sc_hd__or2b_1 _22798_ (.A(_04454_),
    .B_N(_04455_),
    .X(_04466_));
 sky130_fd_sc_hd__o31a_1 _22799_ (.A1(_04268_),
    .A2(_04431_),
    .A3(_04448_),
    .B1(_04452_),
    .X(_04467_));
 sky130_fd_sc_hd__mux2_1 _22800_ (.A0(_04432_),
    .A1(_04431_),
    .S(_04448_),
    .X(_04468_));
 sky130_fd_sc_hd__a21o_1 _22801_ (.A1(_04388_),
    .A2(_04446_),
    .B1(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__nand3_1 _22802_ (.A(_04388_),
    .B(_04446_),
    .C(_04468_),
    .Y(_04470_));
 sky130_fd_sc_hd__and2_1 _22803_ (.A(_04469_),
    .B(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__or2b_1 _22804_ (.A(_04467_),
    .B_N(_04471_),
    .X(_04472_));
 sky130_fd_sc_hd__or2b_1 _22805_ (.A(_04471_),
    .B_N(_04467_),
    .X(_04473_));
 sky130_fd_sc_hd__nand2_1 _22806_ (.A(_04472_),
    .B(_04473_),
    .Y(_04474_));
 sky130_fd_sc_hd__xnor2_1 _22807_ (.A(_04466_),
    .B(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__xnor2_1 _22808_ (.A(_04464_),
    .B(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__or2_1 _22809_ (.A(net666),
    .B(_09804_),
    .X(_04477_));
 sky130_fd_sc_hd__o211a_1 _22810_ (.A1(_09787_),
    .A2(_04476_),
    .B1(_04477_),
    .C1(_03929_),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _22811_ (.A0(\top_inst.deskew_buff_inst.col_input[126] ),
    .A1(_04476_),
    .S(_06140_),
    .X(_04478_));
 sky130_fd_sc_hd__and2_1 _22812_ (.A(_07707_),
    .B(_04478_),
    .X(_04479_));
 sky130_fd_sc_hd__clkbuf_1 _22813_ (.A(_04479_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _22814_ (.A0(_04411_),
    .A1(_04430_),
    .S(_04268_),
    .X(_04480_));
 sky130_fd_sc_hd__xnor2_1 _22815_ (.A(_04444_),
    .B(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__xnor2_1 _22816_ (.A(_04445_),
    .B(_04481_),
    .Y(_04482_));
 sky130_fd_sc_hd__a21oi_2 _22817_ (.A1(_04449_),
    .A2(_04469_),
    .B1(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__and3_1 _22818_ (.A(_04449_),
    .B(_04469_),
    .C(_04482_),
    .X(_04484_));
 sky130_fd_sc_hd__a21o_1 _22819_ (.A1(_04466_),
    .A2(_04462_),
    .B1(_04474_),
    .X(_04485_));
 sky130_fd_sc_hd__o31ai_1 _22820_ (.A1(_04472_),
    .A2(_04483_),
    .A3(_04484_),
    .B1(_04485_),
    .Y(_04486_));
 sky130_fd_sc_hd__a211o_1 _22821_ (.A1(_04364_),
    .A2(_04459_),
    .B1(_04461_),
    .C1(_04486_),
    .X(_04487_));
 sky130_fd_sc_hd__nand2_1 _22822_ (.A(_03700_),
    .B(_03698_),
    .Y(_04488_));
 sky130_fd_sc_hd__a21o_1 _22823_ (.A1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[25] ),
    .A2(_04488_),
    .B1(_03892_),
    .X(_04489_));
 sky130_fd_sc_hd__a31o_1 _22824_ (.A1(_04092_),
    .A2(_04268_),
    .A3(_04489_),
    .B1(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[27] ),
    .X(_04490_));
 sky130_fd_sc_hd__xnor2_1 _22825_ (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[31] ),
    .B(_04483_),
    .Y(_04491_));
 sky130_fd_sc_hd__xnor2_1 _22826_ (.A(_04490_),
    .B(_04491_),
    .Y(_04492_));
 sky130_fd_sc_hd__xnor2_1 _22827_ (.A(_04487_),
    .B(_04492_),
    .Y(_04493_));
 sky130_fd_sc_hd__or2_1 _22828_ (.A(net499),
    .B(_09804_),
    .X(_04494_));
 sky130_fd_sc_hd__o211a_1 _22829_ (.A1(_09787_),
    .A2(_04493_),
    .B1(_04494_),
    .C1(_03929_),
    .X(_00901_));
 sky130_fd_sc_hd__or2_1 _22830_ (.A(\top_inst.skew_buff_inst.row[3].output_reg[0] ),
    .B(_03691_),
    .X(_04495_));
 sky130_fd_sc_hd__o211a_1 _22831_ (.A1(net936),
    .A2(_02877_),
    .B1(_04495_),
    .C1(_03929_),
    .X(_00902_));
 sky130_fd_sc_hd__clkbuf_4 _22832_ (.A(_10583_),
    .X(_04496_));
 sky130_fd_sc_hd__or2_1 _22833_ (.A(\top_inst.skew_buff_inst.row[3].output_reg[1] ),
    .B(_03691_),
    .X(_04497_));
 sky130_fd_sc_hd__buf_2 _22834_ (.A(_02706_),
    .X(_04498_));
 sky130_fd_sc_hd__o211a_1 _22835_ (.A1(net578),
    .A2(_04496_),
    .B1(_04497_),
    .C1(_04498_),
    .X(_00903_));
 sky130_fd_sc_hd__or2_1 _22836_ (.A(\top_inst.skew_buff_inst.row[3].output_reg[2] ),
    .B(_03691_),
    .X(_04499_));
 sky130_fd_sc_hd__o211a_1 _22837_ (.A1(net655),
    .A2(_04496_),
    .B1(_04499_),
    .C1(_04498_),
    .X(_00904_));
 sky130_fd_sc_hd__or2_1 _22838_ (.A(\top_inst.skew_buff_inst.row[3].output_reg[3] ),
    .B(_03691_),
    .X(_04500_));
 sky130_fd_sc_hd__o211a_1 _22839_ (.A1(net406),
    .A2(_04496_),
    .B1(_04500_),
    .C1(_04498_),
    .X(_00905_));
 sky130_fd_sc_hd__or2_1 _22840_ (.A(\top_inst.skew_buff_inst.row[3].output_reg[4] ),
    .B(_03691_),
    .X(_04501_));
 sky130_fd_sc_hd__o211a_1 _22841_ (.A1(net898),
    .A2(_04496_),
    .B1(_04501_),
    .C1(_04498_),
    .X(_00906_));
 sky130_fd_sc_hd__or2_1 _22842_ (.A(\top_inst.skew_buff_inst.row[3].output_reg[5] ),
    .B(_03691_),
    .X(_04502_));
 sky130_fd_sc_hd__o211a_1 _22843_ (.A1(net674),
    .A2(_04496_),
    .B1(_04502_),
    .C1(_04498_),
    .X(_00907_));
 sky130_fd_sc_hd__or2_1 _22844_ (.A(\top_inst.skew_buff_inst.row[3].output_reg[6] ),
    .B(_03691_),
    .X(_04503_));
 sky130_fd_sc_hd__o211a_1 _22845_ (.A1(net394),
    .A2(_04496_),
    .B1(_04503_),
    .C1(_04498_),
    .X(_00908_));
 sky130_fd_sc_hd__buf_2 _22846_ (.A(_06619_),
    .X(_04504_));
 sky130_fd_sc_hd__or2_1 _22847_ (.A(\top_inst.skew_buff_inst.row[3].output_reg[7] ),
    .B(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__o211a_1 _22848_ (.A1(net850),
    .A2(_04496_),
    .B1(_04505_),
    .C1(_04498_),
    .X(_00909_));
 sky130_fd_sc_hd__or2_1 _22849_ (.A(net715),
    .B(_04504_),
    .X(_04506_));
 sky130_fd_sc_hd__o211a_1 _22850_ (.A1(net987),
    .A2(_04496_),
    .B1(_04506_),
    .C1(_04498_),
    .X(_00910_));
 sky130_fd_sc_hd__or2_1 _22851_ (.A(net762),
    .B(_04504_),
    .X(_04507_));
 sky130_fd_sc_hd__o211a_1 _22852_ (.A1(net942),
    .A2(_04496_),
    .B1(_04507_),
    .C1(_04498_),
    .X(_00911_));
 sky130_fd_sc_hd__or2_1 _22853_ (.A(net387),
    .B(_04504_),
    .X(_04508_));
 sky130_fd_sc_hd__o211a_1 _22854_ (.A1(net1039),
    .A2(_04496_),
    .B1(_04508_),
    .C1(_04498_),
    .X(_00912_));
 sky130_fd_sc_hd__clkbuf_4 _22855_ (.A(_10583_),
    .X(_04509_));
 sky130_fd_sc_hd__or2_1 _22856_ (.A(net707),
    .B(_04504_),
    .X(_04510_));
 sky130_fd_sc_hd__clkbuf_4 _22857_ (.A(_02706_),
    .X(_04511_));
 sky130_fd_sc_hd__o211a_1 _22858_ (.A1(net1034),
    .A2(_04509_),
    .B1(_04510_),
    .C1(_04511_),
    .X(_00913_));
 sky130_fd_sc_hd__or2_1 _22859_ (.A(net809),
    .B(_04504_),
    .X(_04512_));
 sky130_fd_sc_hd__o211a_1 _22860_ (.A1(net1043),
    .A2(_04509_),
    .B1(_04512_),
    .C1(_04511_),
    .X(_00914_));
 sky130_fd_sc_hd__or2_1 _22861_ (.A(net828),
    .B(_04504_),
    .X(_04513_));
 sky130_fd_sc_hd__o211a_1 _22862_ (.A1(net986),
    .A2(_04509_),
    .B1(_04513_),
    .C1(_04511_),
    .X(_00915_));
 sky130_fd_sc_hd__or2_1 _22863_ (.A(net294),
    .B(_04504_),
    .X(_04514_));
 sky130_fd_sc_hd__o211a_1 _22864_ (.A1(net1003),
    .A2(_04509_),
    .B1(_04514_),
    .C1(_04511_),
    .X(_00916_));
 sky130_fd_sc_hd__or2_1 _22865_ (.A(net708),
    .B(_04504_),
    .X(_04515_));
 sky130_fd_sc_hd__o211a_1 _22866_ (.A1(net1006),
    .A2(_04509_),
    .B1(_04515_),
    .C1(_04511_),
    .X(_00917_));
 sky130_fd_sc_hd__or2_1 _22867_ (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][0] ),
    .B(_04504_),
    .X(_04516_));
 sky130_fd_sc_hd__o211a_1 _22868_ (.A1(net715),
    .A2(_04509_),
    .B1(_04516_),
    .C1(_04511_),
    .X(_00918_));
 sky130_fd_sc_hd__buf_2 _22869_ (.A(_06619_),
    .X(_04517_));
 sky130_fd_sc_hd__or2_1 _22870_ (.A(net728),
    .B(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__o211a_1 _22871_ (.A1(net762),
    .A2(_04509_),
    .B1(_04518_),
    .C1(_04511_),
    .X(_00919_));
 sky130_fd_sc_hd__or2_1 _22872_ (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][2] ),
    .B(_04517_),
    .X(_04519_));
 sky130_fd_sc_hd__o211a_1 _22873_ (.A1(net387),
    .A2(_04509_),
    .B1(_04519_),
    .C1(_04511_),
    .X(_00920_));
 sky130_fd_sc_hd__or2_1 _22874_ (.A(net296),
    .B(_04517_),
    .X(_04520_));
 sky130_fd_sc_hd__o211a_1 _22875_ (.A1(net707),
    .A2(_04509_),
    .B1(_04520_),
    .C1(_04511_),
    .X(_00921_));
 sky130_fd_sc_hd__or2_1 _22876_ (.A(net784),
    .B(_04517_),
    .X(_04521_));
 sky130_fd_sc_hd__o211a_1 _22877_ (.A1(net809),
    .A2(_04509_),
    .B1(_04521_),
    .C1(_04511_),
    .X(_00922_));
 sky130_fd_sc_hd__clkbuf_4 _22878_ (.A(_10583_),
    .X(_04522_));
 sky130_fd_sc_hd__or2_1 _22879_ (.A(net746),
    .B(_04517_),
    .X(_04523_));
 sky130_fd_sc_hd__buf_2 _22880_ (.A(_02706_),
    .X(_04524_));
 sky130_fd_sc_hd__o211a_1 _22881_ (.A1(net828),
    .A2(_04522_),
    .B1(_04523_),
    .C1(_04524_),
    .X(_00923_));
 sky130_fd_sc_hd__or2_1 _22882_ (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][6] ),
    .B(_04517_),
    .X(_04525_));
 sky130_fd_sc_hd__o211a_1 _22883_ (.A1(net294),
    .A2(_04522_),
    .B1(_04525_),
    .C1(_04524_),
    .X(_00924_));
 sky130_fd_sc_hd__or2_1 _22884_ (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][7] ),
    .B(_04517_),
    .X(_04526_));
 sky130_fd_sc_hd__o211a_1 _22885_ (.A1(net708),
    .A2(_04522_),
    .B1(_04526_),
    .C1(_04524_),
    .X(_00925_));
 sky130_fd_sc_hd__or2_1 _22886_ (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][0] ),
    .B(_04517_),
    .X(_04527_));
 sky130_fd_sc_hd__o211a_1 _22887_ (.A1(net852),
    .A2(_04522_),
    .B1(_04527_),
    .C1(_04524_),
    .X(_00926_));
 sky130_fd_sc_hd__or2_1 _22888_ (.A(net578),
    .B(_04517_),
    .X(_04528_));
 sky130_fd_sc_hd__o211a_1 _22889_ (.A1(net728),
    .A2(_04522_),
    .B1(_04528_),
    .C1(_04524_),
    .X(_00927_));
 sky130_fd_sc_hd__or2_1 _22890_ (.A(net655),
    .B(_04517_),
    .X(_04529_));
 sky130_fd_sc_hd__o211a_1 _22891_ (.A1(net761),
    .A2(_04522_),
    .B1(_04529_),
    .C1(_04524_),
    .X(_00928_));
 sky130_fd_sc_hd__buf_2 _22892_ (.A(_06619_),
    .X(_04530_));
 sky130_fd_sc_hd__or2_1 _22893_ (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][3] ),
    .B(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__o211a_1 _22894_ (.A1(net296),
    .A2(_04522_),
    .B1(_04531_),
    .C1(_04524_),
    .X(_00929_));
 sky130_fd_sc_hd__or2_1 _22895_ (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][4] ),
    .B(_04530_),
    .X(_04532_));
 sky130_fd_sc_hd__o211a_1 _22896_ (.A1(net784),
    .A2(_04522_),
    .B1(_04532_),
    .C1(_04524_),
    .X(_00930_));
 sky130_fd_sc_hd__or2_1 _22897_ (.A(net674),
    .B(_04530_),
    .X(_04533_));
 sky130_fd_sc_hd__o211a_1 _22898_ (.A1(net746),
    .A2(_04522_),
    .B1(_04533_),
    .C1(_04524_),
    .X(_00931_));
 sky130_fd_sc_hd__or2_1 _22899_ (.A(net394),
    .B(_04530_),
    .X(_04534_));
 sky130_fd_sc_hd__o211a_1 _22900_ (.A1(net771),
    .A2(_04522_),
    .B1(_04534_),
    .C1(_04524_),
    .X(_00932_));
 sky130_fd_sc_hd__clkbuf_4 _22901_ (.A(_10583_),
    .X(_04535_));
 sky130_fd_sc_hd__or2_1 _22902_ (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][7] ),
    .B(_04530_),
    .X(_04536_));
 sky130_fd_sc_hd__clkbuf_4 _22903_ (.A(_02706_),
    .X(_04537_));
 sky130_fd_sc_hd__o211a_1 _22904_ (.A1(net764),
    .A2(_04535_),
    .B1(_04536_),
    .C1(_04537_),
    .X(_00933_));
 sky130_fd_sc_hd__or2_1 _22905_ (.A(\top_inst.skew_buff_inst.row[2].output_reg[0] ),
    .B(_04530_),
    .X(_04538_));
 sky130_fd_sc_hd__o211a_1 _22906_ (.A1(net396),
    .A2(_04535_),
    .B1(_04538_),
    .C1(_04537_),
    .X(_00934_));
 sky130_fd_sc_hd__or2_1 _22907_ (.A(\top_inst.skew_buff_inst.row[2].output_reg[1] ),
    .B(_04530_),
    .X(_04539_));
 sky130_fd_sc_hd__o211a_1 _22908_ (.A1(net769),
    .A2(_04535_),
    .B1(_04539_),
    .C1(_04537_),
    .X(_00935_));
 sky130_fd_sc_hd__or2_1 _22909_ (.A(\top_inst.skew_buff_inst.row[2].output_reg[2] ),
    .B(_04530_),
    .X(_04540_));
 sky130_fd_sc_hd__o211a_1 _22910_ (.A1(net766),
    .A2(_04535_),
    .B1(_04540_),
    .C1(_04537_),
    .X(_00936_));
 sky130_fd_sc_hd__or2_1 _22911_ (.A(\top_inst.skew_buff_inst.row[2].output_reg[3] ),
    .B(_04530_),
    .X(_04541_));
 sky130_fd_sc_hd__o211a_1 _22912_ (.A1(net413),
    .A2(_04535_),
    .B1(_04541_),
    .C1(_04537_),
    .X(_00937_));
 sky130_fd_sc_hd__or2_1 _22913_ (.A(\top_inst.skew_buff_inst.row[2].output_reg[4] ),
    .B(_04530_),
    .X(_04542_));
 sky130_fd_sc_hd__o211a_1 _22914_ (.A1(net416),
    .A2(_04535_),
    .B1(_04542_),
    .C1(_04537_),
    .X(_00938_));
 sky130_fd_sc_hd__clkbuf_2 _22915_ (.A(_06619_),
    .X(_04543_));
 sky130_fd_sc_hd__or2_1 _22916_ (.A(\top_inst.skew_buff_inst.row[2].output_reg[5] ),
    .B(_04543_),
    .X(_04544_));
 sky130_fd_sc_hd__o211a_1 _22917_ (.A1(net389),
    .A2(_04535_),
    .B1(_04544_),
    .C1(_04537_),
    .X(_00939_));
 sky130_fd_sc_hd__or2_1 _22918_ (.A(\top_inst.skew_buff_inst.row[2].output_reg[6] ),
    .B(_04543_),
    .X(_04545_));
 sky130_fd_sc_hd__o211a_1 _22919_ (.A1(net380),
    .A2(_04535_),
    .B1(_04545_),
    .C1(_04537_),
    .X(_00940_));
 sky130_fd_sc_hd__or2_1 _22920_ (.A(\top_inst.skew_buff_inst.row[2].output_reg[7] ),
    .B(_04543_),
    .X(_04546_));
 sky130_fd_sc_hd__o211a_1 _22921_ (.A1(net712),
    .A2(_04535_),
    .B1(_04546_),
    .C1(_04537_),
    .X(_00941_));
 sky130_fd_sc_hd__or2_1 _22922_ (.A(net732),
    .B(_04543_),
    .X(_04547_));
 sky130_fd_sc_hd__o211a_1 _22923_ (.A1(net1029),
    .A2(_04535_),
    .B1(_04547_),
    .C1(_04537_),
    .X(_00942_));
 sky130_fd_sc_hd__clkbuf_4 _22924_ (.A(_10583_),
    .X(_04548_));
 sky130_fd_sc_hd__or2_1 _22925_ (.A(net643),
    .B(_04543_),
    .X(_04549_));
 sky130_fd_sc_hd__clkbuf_8 _22926_ (.A(_04868_),
    .X(_04550_));
 sky130_fd_sc_hd__buf_2 _22927_ (.A(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__o211a_1 _22928_ (.A1(net991),
    .A2(_04548_),
    .B1(_04549_),
    .C1(_04551_),
    .X(_00943_));
 sky130_fd_sc_hd__or2_1 _22929_ (.A(net662),
    .B(_04543_),
    .X(_04552_));
 sky130_fd_sc_hd__o211a_1 _22930_ (.A1(net994),
    .A2(_04548_),
    .B1(_04552_),
    .C1(_04551_),
    .X(_00944_));
 sky130_fd_sc_hd__or2_1 _22931_ (.A(net704),
    .B(_04543_),
    .X(_04553_));
 sky130_fd_sc_hd__o211a_1 _22932_ (.A1(net918),
    .A2(_04548_),
    .B1(_04553_),
    .C1(_04551_),
    .X(_00945_));
 sky130_fd_sc_hd__or2_1 _22933_ (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][4] ),
    .B(_04543_),
    .X(_04554_));
 sky130_fd_sc_hd__o211a_1 _22934_ (.A1(net590),
    .A2(_04548_),
    .B1(_04554_),
    .C1(_04551_),
    .X(_00946_));
 sky130_fd_sc_hd__or2_1 _22935_ (.A(net612),
    .B(_04543_),
    .X(_04555_));
 sky130_fd_sc_hd__o211a_1 _22936_ (.A1(net1007),
    .A2(_04548_),
    .B1(_04555_),
    .C1(_04551_),
    .X(_00947_));
 sky130_fd_sc_hd__or2_1 _22937_ (.A(net621),
    .B(_04543_),
    .X(_04556_));
 sky130_fd_sc_hd__o211a_1 _22938_ (.A1(net1037),
    .A2(_04548_),
    .B1(_04556_),
    .C1(_04551_),
    .X(_00948_));
 sky130_fd_sc_hd__buf_2 _22939_ (.A(_04863_),
    .X(_04557_));
 sky130_fd_sc_hd__or2_1 _22940_ (.A(net404),
    .B(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__o211a_1 _22941_ (.A1(net1015),
    .A2(_04548_),
    .B1(_04558_),
    .C1(_04551_),
    .X(_00949_));
 sky130_fd_sc_hd__or2_1 _22942_ (.A(net396),
    .B(_04557_),
    .X(_04559_));
 sky130_fd_sc_hd__o211a_1 _22943_ (.A1(net732),
    .A2(_04548_),
    .B1(_04559_),
    .C1(_04551_),
    .X(_00950_));
 sky130_fd_sc_hd__or2_1 _22944_ (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][1] ),
    .B(_04557_),
    .X(_04560_));
 sky130_fd_sc_hd__o211a_1 _22945_ (.A1(net643),
    .A2(_04548_),
    .B1(_04560_),
    .C1(_04551_),
    .X(_00951_));
 sky130_fd_sc_hd__or2_1 _22946_ (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][2] ),
    .B(_04557_),
    .X(_04561_));
 sky130_fd_sc_hd__o211a_1 _22947_ (.A1(net662),
    .A2(_04548_),
    .B1(_04561_),
    .C1(_04551_),
    .X(_00952_));
 sky130_fd_sc_hd__clkbuf_4 _22948_ (.A(_10583_),
    .X(_04562_));
 sky130_fd_sc_hd__or2_1 _22949_ (.A(net413),
    .B(_04557_),
    .X(_04563_));
 sky130_fd_sc_hd__clkbuf_4 _22950_ (.A(_04550_),
    .X(_04564_));
 sky130_fd_sc_hd__o211a_1 _22951_ (.A1(net704),
    .A2(_04562_),
    .B1(_04563_),
    .C1(_04564_),
    .X(_00953_));
 sky130_fd_sc_hd__or2_1 _22952_ (.A(net416),
    .B(_04557_),
    .X(_04565_));
 sky130_fd_sc_hd__o211a_1 _22953_ (.A1(net681),
    .A2(_04562_),
    .B1(_04565_),
    .C1(_04564_),
    .X(_00954_));
 sky130_fd_sc_hd__or2_1 _22954_ (.A(net389),
    .B(_04557_),
    .X(_04566_));
 sky130_fd_sc_hd__o211a_1 _22955_ (.A1(net612),
    .A2(_04562_),
    .B1(_04566_),
    .C1(_04564_),
    .X(_00955_));
 sky130_fd_sc_hd__or2_1 _22956_ (.A(net380),
    .B(_04557_),
    .X(_04567_));
 sky130_fd_sc_hd__o211a_1 _22957_ (.A1(net621),
    .A2(_04562_),
    .B1(_04567_),
    .C1(_04564_),
    .X(_00956_));
 sky130_fd_sc_hd__or2_1 _22958_ (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][7] ),
    .B(_04557_),
    .X(_04568_));
 sky130_fd_sc_hd__o211a_1 _22959_ (.A1(net404),
    .A2(_04562_),
    .B1(_04568_),
    .C1(_04564_),
    .X(_00957_));
 sky130_fd_sc_hd__or2_1 _22960_ (.A(\top_inst.skew_buff_inst.row[1].output_reg[0] ),
    .B(_04557_),
    .X(_04569_));
 sky130_fd_sc_hd__o211a_1 _22961_ (.A1(net734),
    .A2(_04562_),
    .B1(_04569_),
    .C1(_04564_),
    .X(_00958_));
 sky130_fd_sc_hd__buf_2 _22962_ (.A(_04863_),
    .X(_04570_));
 sky130_fd_sc_hd__or2_1 _22963_ (.A(\top_inst.skew_buff_inst.row[1].output_reg[1] ),
    .B(_04570_),
    .X(_04571_));
 sky130_fd_sc_hd__o211a_1 _22964_ (.A1(net602),
    .A2(_04562_),
    .B1(_04571_),
    .C1(_04564_),
    .X(_00959_));
 sky130_fd_sc_hd__or2_1 _22965_ (.A(\top_inst.skew_buff_inst.row[1].output_reg[2] ),
    .B(_04570_),
    .X(_04572_));
 sky130_fd_sc_hd__o211a_1 _22966_ (.A1(net772),
    .A2(_04562_),
    .B1(_04572_),
    .C1(_04564_),
    .X(_00960_));
 sky130_fd_sc_hd__or2_1 _22967_ (.A(\top_inst.skew_buff_inst.row[1].output_reg[3] ),
    .B(_04570_),
    .X(_04573_));
 sky130_fd_sc_hd__o211a_1 _22968_ (.A1(net702),
    .A2(_04562_),
    .B1(_04573_),
    .C1(_04564_),
    .X(_00961_));
 sky130_fd_sc_hd__or2_1 _22969_ (.A(\top_inst.skew_buff_inst.row[1].output_reg[4] ),
    .B(_04570_),
    .X(_04574_));
 sky130_fd_sc_hd__o211a_1 _22970_ (.A1(net718),
    .A2(_04562_),
    .B1(_04574_),
    .C1(_04564_),
    .X(_00962_));
 sky130_fd_sc_hd__buf_2 _22971_ (.A(_10583_),
    .X(_04575_));
 sky130_fd_sc_hd__or2_1 _22972_ (.A(\top_inst.skew_buff_inst.row[1].output_reg[5] ),
    .B(_04570_),
    .X(_04576_));
 sky130_fd_sc_hd__clkbuf_4 _22973_ (.A(_04550_),
    .X(_04577_));
 sky130_fd_sc_hd__o211a_1 _22974_ (.A1(net881),
    .A2(_04575_),
    .B1(_04576_),
    .C1(_04577_),
    .X(_00963_));
 sky130_fd_sc_hd__or2_1 _22975_ (.A(\top_inst.skew_buff_inst.row[1].output_reg[6] ),
    .B(_04570_),
    .X(_04578_));
 sky130_fd_sc_hd__o211a_1 _22976_ (.A1(net637),
    .A2(_04575_),
    .B1(_04578_),
    .C1(_04577_),
    .X(_00964_));
 sky130_fd_sc_hd__or2_1 _22977_ (.A(\top_inst.skew_buff_inst.row[1].output_reg[7] ),
    .B(_04570_),
    .X(_04579_));
 sky130_fd_sc_hd__o211a_1 _22978_ (.A1(net633),
    .A2(_04575_),
    .B1(_04579_),
    .C1(_04577_),
    .X(_00965_));
 sky130_fd_sc_hd__or2_1 _22979_ (.A(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][0] ),
    .B(_04570_),
    .X(_04580_));
 sky130_fd_sc_hd__o211a_1 _22980_ (.A1(net606),
    .A2(_04575_),
    .B1(_04580_),
    .C1(_04577_),
    .X(_00966_));
 sky130_fd_sc_hd__or2_1 _22981_ (.A(net602),
    .B(_04570_),
    .X(_04581_));
 sky130_fd_sc_hd__o211a_1 _22982_ (.A1(net992),
    .A2(_04575_),
    .B1(_04581_),
    .C1(_04577_),
    .X(_00967_));
 sky130_fd_sc_hd__or2_1 _22983_ (.A(net772),
    .B(_04570_),
    .X(_04582_));
 sky130_fd_sc_hd__o211a_1 _22984_ (.A1(net969),
    .A2(_04575_),
    .B1(_04582_),
    .C1(_04577_),
    .X(_00968_));
 sky130_fd_sc_hd__clkbuf_4 _22985_ (.A(_04863_),
    .X(_04583_));
 sky130_fd_sc_hd__or2_1 _22986_ (.A(net702),
    .B(_04583_),
    .X(_04584_));
 sky130_fd_sc_hd__o211a_1 _22987_ (.A1(net902),
    .A2(_04575_),
    .B1(_04584_),
    .C1(_04577_),
    .X(_00969_));
 sky130_fd_sc_hd__or2_1 _22988_ (.A(net718),
    .B(_04583_),
    .X(_04585_));
 sky130_fd_sc_hd__o211a_1 _22989_ (.A1(net965),
    .A2(_04575_),
    .B1(_04585_),
    .C1(_04577_),
    .X(_00970_));
 sky130_fd_sc_hd__or2_1 _22990_ (.A(net881),
    .B(_04583_),
    .X(_04586_));
 sky130_fd_sc_hd__o211a_1 _22991_ (.A1(net995),
    .A2(_04575_),
    .B1(_04586_),
    .C1(_04577_),
    .X(_00971_));
 sky130_fd_sc_hd__or2_1 _22992_ (.A(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][6] ),
    .B(_04583_),
    .X(_04587_));
 sky130_fd_sc_hd__o211a_1 _22993_ (.A1(net583),
    .A2(_04575_),
    .B1(_04587_),
    .C1(_04577_),
    .X(_00972_));
 sky130_fd_sc_hd__clkbuf_8 _22994_ (.A(_05736_),
    .X(_04588_));
 sky130_fd_sc_hd__or2_1 _22995_ (.A(net633),
    .B(_04583_),
    .X(_04589_));
 sky130_fd_sc_hd__buf_4 _22996_ (.A(_04550_),
    .X(_04590_));
 sky130_fd_sc_hd__o211a_1 _22997_ (.A1(net971),
    .A2(_04588_),
    .B1(_04589_),
    .C1(_04590_),
    .X(_00973_));
 sky130_fd_sc_hd__or2_1 _22998_ (.A(\top_inst.skew_buff_inst.row[0].output_reg[0] ),
    .B(_04583_),
    .X(_04591_));
 sky130_fd_sc_hd__o211a_1 _22999_ (.A1(net903),
    .A2(_04588_),
    .B1(_04591_),
    .C1(_04590_),
    .X(_00974_));
 sky130_fd_sc_hd__or2_1 _23000_ (.A(\top_inst.skew_buff_inst.row[0].output_reg[1] ),
    .B(_04583_),
    .X(_04592_));
 sky130_fd_sc_hd__o211a_1 _23001_ (.A1(net983),
    .A2(_04588_),
    .B1(_04592_),
    .C1(_04590_),
    .X(_00975_));
 sky130_fd_sc_hd__or2_1 _23002_ (.A(\top_inst.skew_buff_inst.row[0].output_reg[2] ),
    .B(_04583_),
    .X(_04593_));
 sky130_fd_sc_hd__o211a_1 _23003_ (.A1(net951),
    .A2(_04588_),
    .B1(_04593_),
    .C1(_04590_),
    .X(_00976_));
 sky130_fd_sc_hd__or2_1 _23004_ (.A(\top_inst.skew_buff_inst.row[0].output_reg[3] ),
    .B(_04583_),
    .X(_04594_));
 sky130_fd_sc_hd__o211a_1 _23005_ (.A1(net979),
    .A2(_04588_),
    .B1(_04594_),
    .C1(_04590_),
    .X(_00977_));
 sky130_fd_sc_hd__or2_1 _23006_ (.A(\top_inst.skew_buff_inst.row[0].output_reg[4] ),
    .B(_04583_),
    .X(_04595_));
 sky130_fd_sc_hd__o211a_1 _23007_ (.A1(net1019),
    .A2(_04588_),
    .B1(_04595_),
    .C1(_04590_),
    .X(_00978_));
 sky130_fd_sc_hd__clkbuf_8 _23008_ (.A(_04863_),
    .X(_04596_));
 sky130_fd_sc_hd__or2_1 _23009_ (.A(\top_inst.skew_buff_inst.row[0].output_reg[5] ),
    .B(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__o211a_1 _23010_ (.A1(net616),
    .A2(_04588_),
    .B1(_04597_),
    .C1(_04590_),
    .X(_00979_));
 sky130_fd_sc_hd__or2_1 _23011_ (.A(net1063),
    .B(_04596_),
    .X(_04598_));
 sky130_fd_sc_hd__o211a_1 _23012_ (.A1(\top_inst.axis_in_inst.inbuf_bus[6] ),
    .A2(_04588_),
    .B1(_04598_),
    .C1(_04590_),
    .X(_00980_));
 sky130_fd_sc_hd__or2_1 _23013_ (.A(\top_inst.skew_buff_inst.row[0].output_reg[7] ),
    .B(_04596_),
    .X(_04599_));
 sky130_fd_sc_hd__o211a_1 _23014_ (.A1(net258),
    .A2(_04588_),
    .B1(_04599_),
    .C1(_04590_),
    .X(_00981_));
 sky130_fd_sc_hd__nand2_2 _23015_ (.A(net33),
    .B(net37),
    .Y(_04600_));
 sky130_fd_sc_hd__buf_4 _23016_ (.A(_04600_),
    .X(_04601_));
 sky130_fd_sc_hd__and2_1 _23017_ (.A(net33),
    .B(net37),
    .X(_04602_));
 sky130_fd_sc_hd__clkbuf_4 _23018_ (.A(_04602_),
    .X(_04603_));
 sky130_fd_sc_hd__or2_1 _23019_ (.A(net903),
    .B(_04603_),
    .X(_04604_));
 sky130_fd_sc_hd__o211a_1 _23020_ (.A1(net1),
    .A2(_04601_),
    .B1(_04604_),
    .C1(_04590_),
    .X(_00982_));
 sky130_fd_sc_hd__or2_1 _23021_ (.A(net983),
    .B(_04603_),
    .X(_04605_));
 sky130_fd_sc_hd__buf_4 _23022_ (.A(_04550_),
    .X(_04606_));
 sky130_fd_sc_hd__o211a_1 _23023_ (.A1(net12),
    .A2(_04601_),
    .B1(_04605_),
    .C1(_04606_),
    .X(_00983_));
 sky130_fd_sc_hd__or2_1 _23024_ (.A(net951),
    .B(_04603_),
    .X(_04607_));
 sky130_fd_sc_hd__o211a_1 _23025_ (.A1(net23),
    .A2(_04601_),
    .B1(_04607_),
    .C1(_04606_),
    .X(_00984_));
 sky130_fd_sc_hd__or2_1 _23026_ (.A(net979),
    .B(_04603_),
    .X(_04608_));
 sky130_fd_sc_hd__o211a_1 _23027_ (.A1(net26),
    .A2(_04601_),
    .B1(_04608_),
    .C1(_04606_),
    .X(_00985_));
 sky130_fd_sc_hd__or2_1 _23028_ (.A(\top_inst.axis_in_inst.inbuf_bus[4] ),
    .B(_04603_),
    .X(_04609_));
 sky130_fd_sc_hd__o211a_1 _23029_ (.A1(net27),
    .A2(_04601_),
    .B1(_04609_),
    .C1(_04606_),
    .X(_00986_));
 sky130_fd_sc_hd__or2_1 _23030_ (.A(net616),
    .B(_04603_),
    .X(_04610_));
 sky130_fd_sc_hd__o211a_1 _23031_ (.A1(net28),
    .A2(_04601_),
    .B1(_04610_),
    .C1(_04606_),
    .X(_00987_));
 sky130_fd_sc_hd__or2_1 _23032_ (.A(\top_inst.axis_in_inst.inbuf_bus[6] ),
    .B(_04603_),
    .X(_04611_));
 sky130_fd_sc_hd__o211a_1 _23033_ (.A1(net29),
    .A2(_04601_),
    .B1(_04611_),
    .C1(_04606_),
    .X(_00988_));
 sky130_fd_sc_hd__or2_1 _23034_ (.A(net1112),
    .B(_04603_),
    .X(_04612_));
 sky130_fd_sc_hd__o211a_1 _23035_ (.A1(net30),
    .A2(_04601_),
    .B1(_04612_),
    .C1(_04606_),
    .X(_00989_));
 sky130_fd_sc_hd__or2_1 _23036_ (.A(net606),
    .B(_04603_),
    .X(_04613_));
 sky130_fd_sc_hd__o211a_1 _23037_ (.A1(net31),
    .A2(_04601_),
    .B1(_04613_),
    .C1(_04606_),
    .X(_00990_));
 sky130_fd_sc_hd__or2_1 _23038_ (.A(\top_inst.axis_in_inst.inbuf_bus[9] ),
    .B(_04603_),
    .X(_04614_));
 sky130_fd_sc_hd__o211a_1 _23039_ (.A1(net32),
    .A2(_04601_),
    .B1(_04614_),
    .C1(_04606_),
    .X(_00991_));
 sky130_fd_sc_hd__clkbuf_4 _23040_ (.A(_04600_),
    .X(_04615_));
 sky130_fd_sc_hd__buf_2 _23041_ (.A(_04602_),
    .X(_04616_));
 sky130_fd_sc_hd__or2_1 _23042_ (.A(net969),
    .B(_04616_),
    .X(_04617_));
 sky130_fd_sc_hd__o211a_1 _23043_ (.A1(net2),
    .A2(_04615_),
    .B1(_04617_),
    .C1(_04606_),
    .X(_00992_));
 sky130_fd_sc_hd__or2_1 _23044_ (.A(net902),
    .B(_04616_),
    .X(_04618_));
 sky130_fd_sc_hd__clkbuf_4 _23045_ (.A(_04550_),
    .X(_04619_));
 sky130_fd_sc_hd__o211a_1 _23046_ (.A1(net3),
    .A2(_04615_),
    .B1(_04618_),
    .C1(_04619_),
    .X(_00993_));
 sky130_fd_sc_hd__or2_1 _23047_ (.A(net965),
    .B(_04616_),
    .X(_04620_));
 sky130_fd_sc_hd__o211a_1 _23048_ (.A1(net4),
    .A2(_04615_),
    .B1(_04620_),
    .C1(_04619_),
    .X(_00994_));
 sky130_fd_sc_hd__or2_1 _23049_ (.A(net995),
    .B(_04616_),
    .X(_04621_));
 sky130_fd_sc_hd__o211a_1 _23050_ (.A1(net5),
    .A2(_04615_),
    .B1(_04621_),
    .C1(_04619_),
    .X(_00995_));
 sky130_fd_sc_hd__or2_1 _23051_ (.A(net583),
    .B(_04616_),
    .X(_04622_));
 sky130_fd_sc_hd__o211a_1 _23052_ (.A1(net6),
    .A2(_04615_),
    .B1(_04622_),
    .C1(_04619_),
    .X(_00996_));
 sky130_fd_sc_hd__or2_1 _23053_ (.A(net971),
    .B(_04616_),
    .X(_04623_));
 sky130_fd_sc_hd__o211a_1 _23054_ (.A1(net7),
    .A2(_04615_),
    .B1(_04623_),
    .C1(_04619_),
    .X(_00997_));
 sky130_fd_sc_hd__or2_1 _23055_ (.A(\top_inst.axis_in_inst.inbuf_bus[16] ),
    .B(_04616_),
    .X(_04624_));
 sky130_fd_sc_hd__o211a_1 _23056_ (.A1(net8),
    .A2(_04615_),
    .B1(_04624_),
    .C1(_04619_),
    .X(_00998_));
 sky130_fd_sc_hd__or2_1 _23057_ (.A(net991),
    .B(_04616_),
    .X(_04625_));
 sky130_fd_sc_hd__o211a_1 _23058_ (.A1(net9),
    .A2(_04615_),
    .B1(_04625_),
    .C1(_04619_),
    .X(_00999_));
 sky130_fd_sc_hd__or2_1 _23059_ (.A(net994),
    .B(_04616_),
    .X(_04626_));
 sky130_fd_sc_hd__o211a_1 _23060_ (.A1(net10),
    .A2(_04615_),
    .B1(_04626_),
    .C1(_04619_),
    .X(_01000_));
 sky130_fd_sc_hd__or2_1 _23061_ (.A(net1111),
    .B(_04616_),
    .X(_04627_));
 sky130_fd_sc_hd__o211a_1 _23062_ (.A1(net11),
    .A2(_04615_),
    .B1(_04627_),
    .C1(_04619_),
    .X(_01001_));
 sky130_fd_sc_hd__clkbuf_4 _23063_ (.A(_04600_),
    .X(_04628_));
 sky130_fd_sc_hd__buf_2 _23064_ (.A(_04602_),
    .X(_04629_));
 sky130_fd_sc_hd__or2_1 _23065_ (.A(net590),
    .B(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__o211a_1 _23066_ (.A1(net13),
    .A2(_04628_),
    .B1(_04630_),
    .C1(_04619_),
    .X(_01002_));
 sky130_fd_sc_hd__or2_1 _23067_ (.A(net1109),
    .B(_04629_),
    .X(_04631_));
 sky130_fd_sc_hd__clkbuf_4 _23068_ (.A(_04550_),
    .X(_04632_));
 sky130_fd_sc_hd__o211a_1 _23069_ (.A1(net14),
    .A2(_04628_),
    .B1(_04631_),
    .C1(_04632_),
    .X(_01003_));
 sky130_fd_sc_hd__or2_1 _23070_ (.A(\top_inst.axis_in_inst.inbuf_bus[22] ),
    .B(_04629_),
    .X(_04633_));
 sky130_fd_sc_hd__o211a_1 _23071_ (.A1(net15),
    .A2(_04628_),
    .B1(_04633_),
    .C1(_04632_),
    .X(_01004_));
 sky130_fd_sc_hd__or2_1 _23072_ (.A(net1110),
    .B(_04629_),
    .X(_04634_));
 sky130_fd_sc_hd__o211a_1 _23073_ (.A1(net16),
    .A2(_04628_),
    .B1(_04634_),
    .C1(_04632_),
    .X(_01005_));
 sky130_fd_sc_hd__or2_1 _23074_ (.A(\top_inst.axis_in_inst.inbuf_bus[24] ),
    .B(_04629_),
    .X(_04635_));
 sky130_fd_sc_hd__o211a_1 _23075_ (.A1(net17),
    .A2(_04628_),
    .B1(_04635_),
    .C1(_04632_),
    .X(_01006_));
 sky130_fd_sc_hd__or2_1 _23076_ (.A(\top_inst.axis_in_inst.inbuf_bus[25] ),
    .B(_04629_),
    .X(_04636_));
 sky130_fd_sc_hd__o211a_1 _23077_ (.A1(net18),
    .A2(_04628_),
    .B1(_04636_),
    .C1(_04632_),
    .X(_01007_));
 sky130_fd_sc_hd__or2_1 _23078_ (.A(\top_inst.axis_in_inst.inbuf_bus[26] ),
    .B(_04629_),
    .X(_04637_));
 sky130_fd_sc_hd__o211a_1 _23079_ (.A1(net19),
    .A2(_04628_),
    .B1(_04637_),
    .C1(_04632_),
    .X(_01008_));
 sky130_fd_sc_hd__or2_1 _23080_ (.A(net1114),
    .B(_04629_),
    .X(_04638_));
 sky130_fd_sc_hd__o211a_1 _23081_ (.A1(net20),
    .A2(_04628_),
    .B1(_04638_),
    .C1(_04632_),
    .X(_01009_));
 sky130_fd_sc_hd__or2_1 _23082_ (.A(\top_inst.axis_in_inst.inbuf_bus[28] ),
    .B(_04629_),
    .X(_04639_));
 sky130_fd_sc_hd__o211a_1 _23083_ (.A1(net21),
    .A2(_04628_),
    .B1(_04639_),
    .C1(_04632_),
    .X(_01010_));
 sky130_fd_sc_hd__or2_1 _23084_ (.A(\top_inst.axis_in_inst.inbuf_bus[29] ),
    .B(_04629_),
    .X(_04640_));
 sky130_fd_sc_hd__o211a_1 _23085_ (.A1(net22),
    .A2(_04628_),
    .B1(_04640_),
    .C1(_04632_),
    .X(_01011_));
 sky130_fd_sc_hd__or2_1 _23086_ (.A(net1115),
    .B(_04602_),
    .X(_04641_));
 sky130_fd_sc_hd__o211a_1 _23087_ (.A1(net24),
    .A2(_04600_),
    .B1(_04641_),
    .C1(_04632_),
    .X(_01012_));
 sky130_fd_sc_hd__or2_1 _23088_ (.A(net1113),
    .B(_04602_),
    .X(_04642_));
 sky130_fd_sc_hd__buf_4 _23089_ (.A(_04550_),
    .X(_04643_));
 sky130_fd_sc_hd__o211a_1 _23090_ (.A1(net25),
    .A2(_04600_),
    .B1(_04642_),
    .C1(_04643_),
    .X(_01013_));
 sky130_fd_sc_hd__inv_2 _23091_ (.A(net33),
    .Y(_04644_));
 sky130_fd_sc_hd__a21oi_1 _23092_ (.A1(_04644_),
    .A2(net37),
    .B1(_04867_),
    .Y(_01014_));
 sky130_fd_sc_hd__nand2_1 _23093_ (.A(net580),
    .B(_10541_),
    .Y(_04645_));
 sky130_fd_sc_hd__a21oi_1 _23094_ (.A1(_09787_),
    .A2(_04645_),
    .B1(_04867_),
    .Y(_01015_));
 sky130_fd_sc_hd__or2_1 _23095_ (.A(net624),
    .B(_05323_),
    .X(_04646_));
 sky130_fd_sc_hd__o211a_1 _23096_ (.A1(net580),
    .A2(_10541_),
    .B1(_04646_),
    .C1(_04643_),
    .X(_01016_));
 sky130_fd_sc_hd__or2_1 _23097_ (.A(net605),
    .B(_05323_),
    .X(_04647_));
 sky130_fd_sc_hd__o211a_1 _23098_ (.A1(net624),
    .A2(_10541_),
    .B1(_04647_),
    .C1(_04643_),
    .X(_01017_));
 sky130_fd_sc_hd__or2_1 _23099_ (.A(net284),
    .B(_05323_),
    .X(_04648_));
 sky130_fd_sc_hd__o211a_1 _23100_ (.A1(net605),
    .A2(_10541_),
    .B1(_04648_),
    .C1(_04643_),
    .X(_01018_));
 sky130_fd_sc_hd__or2_1 _23101_ (.A(\top_inst.valid_pipe[4] ),
    .B(_05323_),
    .X(_04649_));
 sky130_fd_sc_hd__o211a_1 _23102_ (.A1(net284),
    .A2(_10541_),
    .B1(_04649_),
    .C1(_04643_),
    .X(_01019_));
 sky130_fd_sc_hd__or2_1 _23103_ (.A(net354),
    .B(_05323_),
    .X(_04650_));
 sky130_fd_sc_hd__o211a_1 _23104_ (.A1(net653),
    .A2(_10541_),
    .B1(_04650_),
    .C1(_04643_),
    .X(_01020_));
 sky130_fd_sc_hd__or2_1 _23105_ (.A(net331),
    .B(_05323_),
    .X(_04651_));
 sky130_fd_sc_hd__o211a_1 _23106_ (.A1(net354),
    .A2(_10541_),
    .B1(_04651_),
    .C1(_04643_),
    .X(_01021_));
 sky130_fd_sc_hd__or2_1 _23107_ (.A(\top_inst.valid_pipe[7] ),
    .B(_05323_),
    .X(_04652_));
 sky130_fd_sc_hd__o211a_1 _23108_ (.A1(net331),
    .A2(_10541_),
    .B1(_04652_),
    .C1(_04643_),
    .X(_01022_));
 sky130_fd_sc_hd__or2_1 _23109_ (.A(\top_inst.axis_out_inst.out_buff_enabled ),
    .B(_05323_),
    .X(_04653_));
 sky130_fd_sc_hd__o211a_1 _23110_ (.A1(net620),
    .A2(_10541_),
    .B1(_04653_),
    .C1(_04643_),
    .X(_01023_));
 sky130_fd_sc_hd__nand2_1 _23111_ (.A(\top_inst.axis_out_inst.out_buff_enabled ),
    .B(_04857_),
    .Y(_04654_));
 sky130_fd_sc_hd__clkbuf_8 _23112_ (.A(_04654_),
    .X(_04655_));
 sky130_fd_sc_hd__clkbuf_4 _23113_ (.A(_04655_),
    .X(_04656_));
 sky130_fd_sc_hd__and2_1 _23114_ (.A(\top_inst.axis_out_inst.out_buff_enabled ),
    .B(_04857_),
    .X(_04657_));
 sky130_fd_sc_hd__buf_4 _23115_ (.A(_04657_),
    .X(_04658_));
 sky130_fd_sc_hd__buf_2 _23116_ (.A(_04658_),
    .X(_04659_));
 sky130_fd_sc_hd__or2_1 _23117_ (.A(net38),
    .B(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__o211a_1 _23118_ (.A1(net988),
    .A2(_04656_),
    .B1(_04660_),
    .C1(_04643_),
    .X(_01024_));
 sky130_fd_sc_hd__or2_1 _23119_ (.A(net77),
    .B(_04659_),
    .X(_04661_));
 sky130_fd_sc_hd__clkbuf_4 _23120_ (.A(_04550_),
    .X(_04662_));
 sky130_fd_sc_hd__o211a_1 _23121_ (.A1(net787),
    .A2(_04656_),
    .B1(_04661_),
    .C1(_04662_),
    .X(_01025_));
 sky130_fd_sc_hd__or2_1 _23122_ (.A(net88),
    .B(_04659_),
    .X(_04663_));
 sky130_fd_sc_hd__o211a_1 _23123_ (.A1(net677),
    .A2(_04656_),
    .B1(_04663_),
    .C1(_04662_),
    .X(_01026_));
 sky130_fd_sc_hd__or2_1 _23124_ (.A(net99),
    .B(_04659_),
    .X(_04664_));
 sky130_fd_sc_hd__o211a_1 _23125_ (.A1(net463),
    .A2(_04656_),
    .B1(_04664_),
    .C1(_04662_),
    .X(_01027_));
 sky130_fd_sc_hd__or2_1 _23126_ (.A(net110),
    .B(_04659_),
    .X(_04665_));
 sky130_fd_sc_hd__o211a_1 _23127_ (.A1(net422),
    .A2(_04656_),
    .B1(_04665_),
    .C1(_04662_),
    .X(_01028_));
 sky130_fd_sc_hd__or2_1 _23128_ (.A(net121),
    .B(_04659_),
    .X(_04666_));
 sky130_fd_sc_hd__o211a_1 _23129_ (.A1(net686),
    .A2(_04656_),
    .B1(_04666_),
    .C1(_04662_),
    .X(_01029_));
 sky130_fd_sc_hd__or2_1 _23130_ (.A(net132),
    .B(_04659_),
    .X(_04667_));
 sky130_fd_sc_hd__o211a_1 _23131_ (.A1(net541),
    .A2(_04656_),
    .B1(_04667_),
    .C1(_04662_),
    .X(_01030_));
 sky130_fd_sc_hd__or2_1 _23132_ (.A(net143),
    .B(_04659_),
    .X(_04668_));
 sky130_fd_sc_hd__o211a_1 _23133_ (.A1(net755),
    .A2(_04656_),
    .B1(_04668_),
    .C1(_04662_),
    .X(_01031_));
 sky130_fd_sc_hd__or2_1 _23134_ (.A(net154),
    .B(_04659_),
    .X(_04669_));
 sky130_fd_sc_hd__o211a_1 _23135_ (.A1(net310),
    .A2(_04656_),
    .B1(_04669_),
    .C1(_04662_),
    .X(_01032_));
 sky130_fd_sc_hd__or2_1 _23136_ (.A(net165),
    .B(_04659_),
    .X(_04670_));
 sky130_fd_sc_hd__o211a_1 _23137_ (.A1(net661),
    .A2(_04656_),
    .B1(_04670_),
    .C1(_04662_),
    .X(_01033_));
 sky130_fd_sc_hd__clkbuf_4 _23138_ (.A(_04655_),
    .X(_04671_));
 sky130_fd_sc_hd__buf_2 _23139_ (.A(_04658_),
    .X(_04672_));
 sky130_fd_sc_hd__or2_1 _23140_ (.A(net49),
    .B(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__o211a_1 _23141_ (.A1(net440),
    .A2(_04671_),
    .B1(_04673_),
    .C1(_04662_),
    .X(_01034_));
 sky130_fd_sc_hd__or2_1 _23142_ (.A(net60),
    .B(_04672_),
    .X(_04674_));
 sky130_fd_sc_hd__clkbuf_4 _23143_ (.A(_04550_),
    .X(_04675_));
 sky130_fd_sc_hd__o211a_1 _23144_ (.A1(net632),
    .A2(_04671_),
    .B1(_04674_),
    .C1(_04675_),
    .X(_01035_));
 sky130_fd_sc_hd__or2_1 _23145_ (.A(net69),
    .B(_04672_),
    .X(_04676_));
 sky130_fd_sc_hd__o211a_1 _23146_ (.A1(net618),
    .A2(_04671_),
    .B1(_04676_),
    .C1(_04675_),
    .X(_01036_));
 sky130_fd_sc_hd__or2_1 _23147_ (.A(net70),
    .B(_04672_),
    .X(_04677_));
 sky130_fd_sc_hd__o211a_1 _23148_ (.A1(net317),
    .A2(_04671_),
    .B1(_04677_),
    .C1(_04675_),
    .X(_01037_));
 sky130_fd_sc_hd__or2_1 _23149_ (.A(net71),
    .B(_04672_),
    .X(_04678_));
 sky130_fd_sc_hd__o211a_1 _23150_ (.A1(net359),
    .A2(_04671_),
    .B1(_04678_),
    .C1(_04675_),
    .X(_01038_));
 sky130_fd_sc_hd__or2_1 _23151_ (.A(net72),
    .B(_04672_),
    .X(_04679_));
 sky130_fd_sc_hd__o211a_1 _23152_ (.A1(net955),
    .A2(_04671_),
    .B1(_04679_),
    .C1(_04675_),
    .X(_01039_));
 sky130_fd_sc_hd__or2_1 _23153_ (.A(net73),
    .B(_04672_),
    .X(_04680_));
 sky130_fd_sc_hd__o211a_1 _23154_ (.A1(net832),
    .A2(_04671_),
    .B1(_04680_),
    .C1(_04675_),
    .X(_01040_));
 sky130_fd_sc_hd__or2_1 _23155_ (.A(net74),
    .B(_04672_),
    .X(_04681_));
 sky130_fd_sc_hd__o211a_1 _23156_ (.A1(net485),
    .A2(_04671_),
    .B1(_04681_),
    .C1(_04675_),
    .X(_01041_));
 sky130_fd_sc_hd__or2_1 _23157_ (.A(net75),
    .B(_04672_),
    .X(_04682_));
 sky130_fd_sc_hd__o211a_1 _23158_ (.A1(net774),
    .A2(_04671_),
    .B1(_04682_),
    .C1(_04675_),
    .X(_01042_));
 sky130_fd_sc_hd__or2_1 _23159_ (.A(net76),
    .B(_04672_),
    .X(_04683_));
 sky130_fd_sc_hd__o211a_1 _23160_ (.A1(net830),
    .A2(_04671_),
    .B1(_04683_),
    .C1(_04675_),
    .X(_01043_));
 sky130_fd_sc_hd__clkbuf_8 _23161_ (.A(_04654_),
    .X(_04684_));
 sky130_fd_sc_hd__clkbuf_4 _23162_ (.A(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__clkbuf_8 _23163_ (.A(_04657_),
    .X(_04686_));
 sky130_fd_sc_hd__buf_2 _23164_ (.A(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__or2_1 _23165_ (.A(net78),
    .B(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__o211a_1 _23166_ (.A1(net382),
    .A2(_04685_),
    .B1(_04688_),
    .C1(_04675_),
    .X(_01044_));
 sky130_fd_sc_hd__or2_1 _23167_ (.A(net79),
    .B(_04687_),
    .X(_04689_));
 sky130_fd_sc_hd__clkbuf_8 _23168_ (.A(_04868_),
    .X(_04690_));
 sky130_fd_sc_hd__clkbuf_4 _23169_ (.A(_04690_),
    .X(_04691_));
 sky130_fd_sc_hd__o211a_1 _23170_ (.A1(net799),
    .A2(_04685_),
    .B1(_04689_),
    .C1(_04691_),
    .X(_01045_));
 sky130_fd_sc_hd__or2_1 _23171_ (.A(net80),
    .B(_04687_),
    .X(_04692_));
 sky130_fd_sc_hd__o211a_1 _23172_ (.A1(net870),
    .A2(_04685_),
    .B1(_04692_),
    .C1(_04691_),
    .X(_01046_));
 sky130_fd_sc_hd__or2_1 _23173_ (.A(net81),
    .B(_04687_),
    .X(_04693_));
 sky130_fd_sc_hd__o211a_1 _23174_ (.A1(net843),
    .A2(_04685_),
    .B1(_04693_),
    .C1(_04691_),
    .X(_01047_));
 sky130_fd_sc_hd__or2_1 _23175_ (.A(net82),
    .B(_04687_),
    .X(_04694_));
 sky130_fd_sc_hd__o211a_1 _23176_ (.A1(net379),
    .A2(_04685_),
    .B1(_04694_),
    .C1(_04691_),
    .X(_01048_));
 sky130_fd_sc_hd__or2_1 _23177_ (.A(net83),
    .B(_04687_),
    .X(_04695_));
 sky130_fd_sc_hd__o211a_1 _23178_ (.A1(net548),
    .A2(_04685_),
    .B1(_04695_),
    .C1(_04691_),
    .X(_01049_));
 sky130_fd_sc_hd__or2_1 _23179_ (.A(net84),
    .B(_04687_),
    .X(_04696_));
 sky130_fd_sc_hd__o211a_1 _23180_ (.A1(net723),
    .A2(_04685_),
    .B1(_04696_),
    .C1(_04691_),
    .X(_01050_));
 sky130_fd_sc_hd__or2_1 _23181_ (.A(net85),
    .B(_04687_),
    .X(_04697_));
 sky130_fd_sc_hd__o211a_1 _23182_ (.A1(net768),
    .A2(_04685_),
    .B1(_04697_),
    .C1(_04691_),
    .X(_01051_));
 sky130_fd_sc_hd__or2_1 _23183_ (.A(net86),
    .B(_04687_),
    .X(_04698_));
 sky130_fd_sc_hd__o211a_1 _23184_ (.A1(net749),
    .A2(_04685_),
    .B1(_04698_),
    .C1(_04691_),
    .X(_01052_));
 sky130_fd_sc_hd__or2_1 _23185_ (.A(net87),
    .B(_04687_),
    .X(_04699_));
 sky130_fd_sc_hd__o211a_1 _23186_ (.A1(net736),
    .A2(_04685_),
    .B1(_04699_),
    .C1(_04691_),
    .X(_01053_));
 sky130_fd_sc_hd__clkbuf_4 _23187_ (.A(_04684_),
    .X(_04700_));
 sky130_fd_sc_hd__buf_2 _23188_ (.A(_04686_),
    .X(_04701_));
 sky130_fd_sc_hd__or2_1 _23189_ (.A(net89),
    .B(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__o211a_1 _23190_ (.A1(net492),
    .A2(_04700_),
    .B1(_04702_),
    .C1(_04691_),
    .X(_01054_));
 sky130_fd_sc_hd__or2_1 _23191_ (.A(net90),
    .B(_04701_),
    .X(_04703_));
 sky130_fd_sc_hd__clkbuf_4 _23192_ (.A(_04690_),
    .X(_04704_));
 sky130_fd_sc_hd__o211a_1 _23193_ (.A1(net972),
    .A2(_04700_),
    .B1(_04703_),
    .C1(_04704_),
    .X(_01055_));
 sky130_fd_sc_hd__or2_1 _23194_ (.A(net91),
    .B(_04701_),
    .X(_04705_));
 sky130_fd_sc_hd__o211a_1 _23195_ (.A1(net493),
    .A2(_04700_),
    .B1(_04705_),
    .C1(_04704_),
    .X(_01056_));
 sky130_fd_sc_hd__or2_1 _23196_ (.A(net92),
    .B(_04701_),
    .X(_04706_));
 sky130_fd_sc_hd__o211a_1 _23197_ (.A1(net673),
    .A2(_04700_),
    .B1(_04706_),
    .C1(_04704_),
    .X(_01057_));
 sky130_fd_sc_hd__or2_1 _23198_ (.A(net93),
    .B(_04701_),
    .X(_04707_));
 sky130_fd_sc_hd__o211a_1 _23199_ (.A1(net789),
    .A2(_04700_),
    .B1(_04707_),
    .C1(_04704_),
    .X(_01058_));
 sky130_fd_sc_hd__or2_1 _23200_ (.A(net94),
    .B(_04701_),
    .X(_04708_));
 sky130_fd_sc_hd__o211a_1 _23201_ (.A1(net844),
    .A2(_04700_),
    .B1(_04708_),
    .C1(_04704_),
    .X(_01059_));
 sky130_fd_sc_hd__or2_1 _23202_ (.A(net95),
    .B(_04701_),
    .X(_04709_));
 sky130_fd_sc_hd__o211a_1 _23203_ (.A1(net378),
    .A2(_04700_),
    .B1(_04709_),
    .C1(_04704_),
    .X(_01060_));
 sky130_fd_sc_hd__or2_1 _23204_ (.A(net96),
    .B(_04701_),
    .X(_04710_));
 sky130_fd_sc_hd__o211a_1 _23205_ (.A1(net676),
    .A2(_04700_),
    .B1(_04710_),
    .C1(_04704_),
    .X(_01061_));
 sky130_fd_sc_hd__or2_1 _23206_ (.A(net97),
    .B(_04701_),
    .X(_04711_));
 sky130_fd_sc_hd__o211a_1 _23207_ (.A1(net845),
    .A2(_04700_),
    .B1(_04711_),
    .C1(_04704_),
    .X(_01062_));
 sky130_fd_sc_hd__or2_1 _23208_ (.A(net98),
    .B(_04701_),
    .X(_04712_));
 sky130_fd_sc_hd__o211a_1 _23209_ (.A1(net665),
    .A2(_04700_),
    .B1(_04712_),
    .C1(_04704_),
    .X(_01063_));
 sky130_fd_sc_hd__clkbuf_4 _23210_ (.A(_04684_),
    .X(_04713_));
 sky130_fd_sc_hd__buf_2 _23211_ (.A(_04686_),
    .X(_04714_));
 sky130_fd_sc_hd__or2_1 _23212_ (.A(net100),
    .B(_04714_),
    .X(_04715_));
 sky130_fd_sc_hd__o211a_1 _23213_ (.A1(net595),
    .A2(_04713_),
    .B1(_04715_),
    .C1(_04704_),
    .X(_01064_));
 sky130_fd_sc_hd__or2_1 _23214_ (.A(net101),
    .B(_04714_),
    .X(_04716_));
 sky130_fd_sc_hd__clkbuf_4 _23215_ (.A(_04690_),
    .X(_04717_));
 sky130_fd_sc_hd__o211a_1 _23216_ (.A1(net822),
    .A2(_04713_),
    .B1(_04716_),
    .C1(_04717_),
    .X(_01065_));
 sky130_fd_sc_hd__or2_1 _23217_ (.A(net102),
    .B(_04714_),
    .X(_04718_));
 sky130_fd_sc_hd__o211a_1 _23218_ (.A1(net613),
    .A2(_04713_),
    .B1(_04718_),
    .C1(_04717_),
    .X(_01066_));
 sky130_fd_sc_hd__or2_1 _23219_ (.A(net103),
    .B(_04714_),
    .X(_04719_));
 sky130_fd_sc_hd__o211a_1 _23220_ (.A1(net610),
    .A2(_04713_),
    .B1(_04719_),
    .C1(_04717_),
    .X(_01067_));
 sky130_fd_sc_hd__or2_1 _23221_ (.A(net104),
    .B(_04714_),
    .X(_04720_));
 sky130_fd_sc_hd__o211a_1 _23222_ (.A1(net513),
    .A2(_04713_),
    .B1(_04720_),
    .C1(_04717_),
    .X(_01068_));
 sky130_fd_sc_hd__or2_1 _23223_ (.A(net105),
    .B(_04714_),
    .X(_04721_));
 sky130_fd_sc_hd__o211a_1 _23224_ (.A1(net763),
    .A2(_04713_),
    .B1(_04721_),
    .C1(_04717_),
    .X(_01069_));
 sky130_fd_sc_hd__or2_1 _23225_ (.A(net106),
    .B(_04714_),
    .X(_04722_));
 sky130_fd_sc_hd__o211a_1 _23226_ (.A1(net731),
    .A2(_04713_),
    .B1(_04722_),
    .C1(_04717_),
    .X(_01070_));
 sky130_fd_sc_hd__or2_1 _23227_ (.A(net107),
    .B(_04714_),
    .X(_04723_));
 sky130_fd_sc_hd__o211a_1 _23228_ (.A1(net651),
    .A2(_04713_),
    .B1(_04723_),
    .C1(_04717_),
    .X(_01071_));
 sky130_fd_sc_hd__or2_1 _23229_ (.A(net108),
    .B(_04714_),
    .X(_04724_));
 sky130_fd_sc_hd__o211a_1 _23230_ (.A1(net553),
    .A2(_04713_),
    .B1(_04724_),
    .C1(_04717_),
    .X(_01072_));
 sky130_fd_sc_hd__or2_1 _23231_ (.A(net109),
    .B(_04714_),
    .X(_04725_));
 sky130_fd_sc_hd__o211a_1 _23232_ (.A1(net699),
    .A2(_04713_),
    .B1(_04725_),
    .C1(_04717_),
    .X(_01073_));
 sky130_fd_sc_hd__clkbuf_4 _23233_ (.A(_04684_),
    .X(_04726_));
 sky130_fd_sc_hd__clkbuf_4 _23234_ (.A(_04686_),
    .X(_04727_));
 sky130_fd_sc_hd__or2_1 _23235_ (.A(net111),
    .B(_04727_),
    .X(_04728_));
 sky130_fd_sc_hd__o211a_1 _23236_ (.A1(net796),
    .A2(_04726_),
    .B1(_04728_),
    .C1(_04717_),
    .X(_01074_));
 sky130_fd_sc_hd__or2_1 _23237_ (.A(net112),
    .B(_04727_),
    .X(_04729_));
 sky130_fd_sc_hd__clkbuf_4 _23238_ (.A(_04690_),
    .X(_04730_));
 sky130_fd_sc_hd__o211a_1 _23239_ (.A1(net693),
    .A2(_04726_),
    .B1(_04729_),
    .C1(_04730_),
    .X(_01075_));
 sky130_fd_sc_hd__or2_1 _23240_ (.A(net113),
    .B(_04727_),
    .X(_04731_));
 sky130_fd_sc_hd__o211a_1 _23241_ (.A1(net978),
    .A2(_04726_),
    .B1(_04731_),
    .C1(_04730_),
    .X(_01076_));
 sky130_fd_sc_hd__or2_1 _23242_ (.A(net114),
    .B(_04727_),
    .X(_04732_));
 sky130_fd_sc_hd__o211a_1 _23243_ (.A1(net873),
    .A2(_04726_),
    .B1(_04732_),
    .C1(_04730_),
    .X(_01077_));
 sky130_fd_sc_hd__or2_1 _23244_ (.A(net115),
    .B(_04727_),
    .X(_04733_));
 sky130_fd_sc_hd__o211a_1 _23245_ (.A1(net802),
    .A2(_04726_),
    .B1(_04733_),
    .C1(_04730_),
    .X(_01078_));
 sky130_fd_sc_hd__or2_1 _23246_ (.A(net116),
    .B(_04727_),
    .X(_04734_));
 sky130_fd_sc_hd__o211a_1 _23247_ (.A1(net945),
    .A2(_04726_),
    .B1(_04734_),
    .C1(_04730_),
    .X(_01079_));
 sky130_fd_sc_hd__or2_1 _23248_ (.A(net117),
    .B(_04727_),
    .X(_04735_));
 sky130_fd_sc_hd__o211a_1 _23249_ (.A1(net838),
    .A2(_04726_),
    .B1(_04735_),
    .C1(_04730_),
    .X(_01080_));
 sky130_fd_sc_hd__or2_1 _23250_ (.A(net118),
    .B(_04727_),
    .X(_04736_));
 sky130_fd_sc_hd__o211a_1 _23251_ (.A1(net821),
    .A2(_04726_),
    .B1(_04736_),
    .C1(_04730_),
    .X(_01081_));
 sky130_fd_sc_hd__or2_1 _23252_ (.A(net119),
    .B(_04727_),
    .X(_04737_));
 sky130_fd_sc_hd__o211a_1 _23253_ (.A1(net1025),
    .A2(_04726_),
    .B1(_04737_),
    .C1(_04730_),
    .X(_01082_));
 sky130_fd_sc_hd__or2_1 _23254_ (.A(net120),
    .B(_04727_),
    .X(_04738_));
 sky130_fd_sc_hd__o211a_1 _23255_ (.A1(net920),
    .A2(_04726_),
    .B1(_04738_),
    .C1(_04730_),
    .X(_01083_));
 sky130_fd_sc_hd__buf_4 _23256_ (.A(_04684_),
    .X(_04739_));
 sky130_fd_sc_hd__clkbuf_4 _23257_ (.A(_04686_),
    .X(_04740_));
 sky130_fd_sc_hd__or2_1 _23258_ (.A(net122),
    .B(_04740_),
    .X(_04741_));
 sky130_fd_sc_hd__o211a_1 _23259_ (.A1(net752),
    .A2(_04739_),
    .B1(_04741_),
    .C1(_04730_),
    .X(_01084_));
 sky130_fd_sc_hd__or2_1 _23260_ (.A(net123),
    .B(_04740_),
    .X(_04742_));
 sky130_fd_sc_hd__buf_4 _23261_ (.A(_04690_),
    .X(_04743_));
 sky130_fd_sc_hd__o211a_1 _23262_ (.A1(net1059),
    .A2(_04739_),
    .B1(_04742_),
    .C1(_04743_),
    .X(_01085_));
 sky130_fd_sc_hd__or2_1 _23263_ (.A(net124),
    .B(_04740_),
    .X(_04744_));
 sky130_fd_sc_hd__o211a_1 _23264_ (.A1(net730),
    .A2(_04739_),
    .B1(_04744_),
    .C1(_04743_),
    .X(_01086_));
 sky130_fd_sc_hd__or2_1 _23265_ (.A(net125),
    .B(_04740_),
    .X(_04745_));
 sky130_fd_sc_hd__o211a_1 _23266_ (.A1(net1023),
    .A2(_04739_),
    .B1(_04745_),
    .C1(_04743_),
    .X(_01087_));
 sky130_fd_sc_hd__or2_1 _23267_ (.A(net126),
    .B(_04740_),
    .X(_04746_));
 sky130_fd_sc_hd__o211a_1 _23268_ (.A1(net776),
    .A2(_04739_),
    .B1(_04746_),
    .C1(_04743_),
    .X(_01088_));
 sky130_fd_sc_hd__or2_1 _23269_ (.A(net127),
    .B(_04740_),
    .X(_04747_));
 sky130_fd_sc_hd__o211a_1 _23270_ (.A1(net622),
    .A2(_04739_),
    .B1(_04747_),
    .C1(_04743_),
    .X(_01089_));
 sky130_fd_sc_hd__or2_1 _23271_ (.A(net128),
    .B(_04740_),
    .X(_04748_));
 sky130_fd_sc_hd__o211a_1 _23272_ (.A1(net364),
    .A2(_04739_),
    .B1(_04748_),
    .C1(_04743_),
    .X(_01090_));
 sky130_fd_sc_hd__or2_1 _23273_ (.A(net129),
    .B(_04740_),
    .X(_04749_));
 sky130_fd_sc_hd__o211a_1 _23274_ (.A1(net377),
    .A2(_04739_),
    .B1(_04749_),
    .C1(_04743_),
    .X(_01091_));
 sky130_fd_sc_hd__or2_1 _23275_ (.A(net130),
    .B(_04740_),
    .X(_04750_));
 sky130_fd_sc_hd__o211a_1 _23276_ (.A1(net940),
    .A2(_04739_),
    .B1(_04750_),
    .C1(_04743_),
    .X(_01092_));
 sky130_fd_sc_hd__or2_1 _23277_ (.A(net131),
    .B(_04740_),
    .X(_04751_));
 sky130_fd_sc_hd__o211a_1 _23278_ (.A1(net690),
    .A2(_04739_),
    .B1(_04751_),
    .C1(_04743_),
    .X(_01093_));
 sky130_fd_sc_hd__clkbuf_4 _23279_ (.A(_04684_),
    .X(_04752_));
 sky130_fd_sc_hd__clkbuf_2 _23280_ (.A(_04686_),
    .X(_04753_));
 sky130_fd_sc_hd__or2_1 _23281_ (.A(net133),
    .B(_04753_),
    .X(_04754_));
 sky130_fd_sc_hd__o211a_1 _23282_ (.A1(net476),
    .A2(_04752_),
    .B1(_04754_),
    .C1(_04743_),
    .X(_01094_));
 sky130_fd_sc_hd__or2_1 _23283_ (.A(net134),
    .B(_04753_),
    .X(_04755_));
 sky130_fd_sc_hd__clkbuf_4 _23284_ (.A(_04690_),
    .X(_04756_));
 sky130_fd_sc_hd__o211a_1 _23285_ (.A1(net489),
    .A2(_04752_),
    .B1(_04755_),
    .C1(_04756_),
    .X(_01095_));
 sky130_fd_sc_hd__or2_1 _23286_ (.A(net135),
    .B(_04753_),
    .X(_04757_));
 sky130_fd_sc_hd__o211a_1 _23287_ (.A1(net757),
    .A2(_04752_),
    .B1(_04757_),
    .C1(_04756_),
    .X(_01096_));
 sky130_fd_sc_hd__or2_1 _23288_ (.A(net136),
    .B(_04753_),
    .X(_04758_));
 sky130_fd_sc_hd__o211a_1 _23289_ (.A1(net645),
    .A2(_04752_),
    .B1(_04758_),
    .C1(_04756_),
    .X(_01097_));
 sky130_fd_sc_hd__or2_1 _23290_ (.A(net137),
    .B(_04753_),
    .X(_04759_));
 sky130_fd_sc_hd__o211a_1 _23291_ (.A1(net743),
    .A2(_04752_),
    .B1(_04759_),
    .C1(_04756_),
    .X(_01098_));
 sky130_fd_sc_hd__or2_1 _23292_ (.A(net138),
    .B(_04753_),
    .X(_04760_));
 sky130_fd_sc_hd__o211a_1 _23293_ (.A1(net727),
    .A2(_04752_),
    .B1(_04760_),
    .C1(_04756_),
    .X(_01099_));
 sky130_fd_sc_hd__or2_1 _23294_ (.A(net139),
    .B(_04753_),
    .X(_04761_));
 sky130_fd_sc_hd__o211a_1 _23295_ (.A1(net705),
    .A2(_04752_),
    .B1(_04761_),
    .C1(_04756_),
    .X(_01100_));
 sky130_fd_sc_hd__or2_1 _23296_ (.A(net140),
    .B(_04753_),
    .X(_04762_));
 sky130_fd_sc_hd__o211a_1 _23297_ (.A1(net468),
    .A2(_04752_),
    .B1(_04762_),
    .C1(_04756_),
    .X(_01101_));
 sky130_fd_sc_hd__or2_1 _23298_ (.A(net141),
    .B(_04753_),
    .X(_04763_));
 sky130_fd_sc_hd__o211a_1 _23299_ (.A1(net804),
    .A2(_04752_),
    .B1(_04763_),
    .C1(_04756_),
    .X(_01102_));
 sky130_fd_sc_hd__or2_1 _23300_ (.A(net142),
    .B(_04753_),
    .X(_04764_));
 sky130_fd_sc_hd__o211a_1 _23301_ (.A1(net687),
    .A2(_04752_),
    .B1(_04764_),
    .C1(_04756_),
    .X(_01103_));
 sky130_fd_sc_hd__clkbuf_4 _23302_ (.A(_04684_),
    .X(_04765_));
 sky130_fd_sc_hd__buf_2 _23303_ (.A(_04686_),
    .X(_04766_));
 sky130_fd_sc_hd__or2_1 _23304_ (.A(net144),
    .B(_04766_),
    .X(_04767_));
 sky130_fd_sc_hd__o211a_1 _23305_ (.A1(net927),
    .A2(_04765_),
    .B1(_04767_),
    .C1(_04756_),
    .X(_01104_));
 sky130_fd_sc_hd__or2_1 _23306_ (.A(net145),
    .B(_04766_),
    .X(_04768_));
 sky130_fd_sc_hd__clkbuf_4 _23307_ (.A(_04690_),
    .X(_04769_));
 sky130_fd_sc_hd__o211a_1 _23308_ (.A1(net462),
    .A2(_04765_),
    .B1(_04768_),
    .C1(_04769_),
    .X(_01105_));
 sky130_fd_sc_hd__or2_1 _23309_ (.A(net146),
    .B(_04766_),
    .X(_04770_));
 sky130_fd_sc_hd__o211a_1 _23310_ (.A1(net537),
    .A2(_04765_),
    .B1(_04770_),
    .C1(_04769_),
    .X(_01106_));
 sky130_fd_sc_hd__or2_1 _23311_ (.A(net147),
    .B(_04766_),
    .X(_04771_));
 sky130_fd_sc_hd__o211a_1 _23312_ (.A1(net742),
    .A2(_04765_),
    .B1(_04771_),
    .C1(_04769_),
    .X(_01107_));
 sky130_fd_sc_hd__or2_1 _23313_ (.A(net148),
    .B(_04766_),
    .X(_04772_));
 sky130_fd_sc_hd__o211a_1 _23314_ (.A1(net393),
    .A2(_04765_),
    .B1(_04772_),
    .C1(_04769_),
    .X(_01108_));
 sky130_fd_sc_hd__or2_1 _23315_ (.A(net149),
    .B(_04766_),
    .X(_04773_));
 sky130_fd_sc_hd__o211a_1 _23316_ (.A1(net391),
    .A2(_04765_),
    .B1(_04773_),
    .C1(_04769_),
    .X(_01109_));
 sky130_fd_sc_hd__or2_1 _23317_ (.A(net150),
    .B(_04766_),
    .X(_04774_));
 sky130_fd_sc_hd__o211a_1 _23318_ (.A1(net658),
    .A2(_04765_),
    .B1(_04774_),
    .C1(_04769_),
    .X(_01110_));
 sky130_fd_sc_hd__or2_1 _23319_ (.A(net151),
    .B(_04766_),
    .X(_04775_));
 sky130_fd_sc_hd__o211a_1 _23320_ (.A1(net629),
    .A2(_04765_),
    .B1(_04775_),
    .C1(_04769_),
    .X(_01111_));
 sky130_fd_sc_hd__or2_1 _23321_ (.A(net152),
    .B(_04766_),
    .X(_04776_));
 sky130_fd_sc_hd__o211a_1 _23322_ (.A1(net657),
    .A2(_04765_),
    .B1(_04776_),
    .C1(_04769_),
    .X(_01112_));
 sky130_fd_sc_hd__or2_1 _23323_ (.A(net153),
    .B(_04766_),
    .X(_04777_));
 sky130_fd_sc_hd__o211a_1 _23324_ (.A1(net415),
    .A2(_04765_),
    .B1(_04777_),
    .C1(_04769_),
    .X(_01113_));
 sky130_fd_sc_hd__buf_4 _23325_ (.A(_04684_),
    .X(_04778_));
 sky130_fd_sc_hd__buf_4 _23326_ (.A(_04686_),
    .X(_04779_));
 sky130_fd_sc_hd__or2_1 _23327_ (.A(net155),
    .B(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__o211a_1 _23328_ (.A1(net694),
    .A2(_04778_),
    .B1(_04780_),
    .C1(_04769_),
    .X(_01114_));
 sky130_fd_sc_hd__or2_1 _23329_ (.A(net156),
    .B(_04779_),
    .X(_04781_));
 sky130_fd_sc_hd__buf_4 _23330_ (.A(_04690_),
    .X(_04782_));
 sky130_fd_sc_hd__o211a_1 _23331_ (.A1(net599),
    .A2(_04778_),
    .B1(_04781_),
    .C1(_04782_),
    .X(_01115_));
 sky130_fd_sc_hd__or2_1 _23332_ (.A(net157),
    .B(_04779_),
    .X(_04783_));
 sky130_fd_sc_hd__o211a_1 _23333_ (.A1(net434),
    .A2(_04778_),
    .B1(_04783_),
    .C1(_04782_),
    .X(_01116_));
 sky130_fd_sc_hd__or2_1 _23334_ (.A(net158),
    .B(_04779_),
    .X(_04784_));
 sky130_fd_sc_hd__o211a_1 _23335_ (.A1(net831),
    .A2(_04778_),
    .B1(_04784_),
    .C1(_04782_),
    .X(_01117_));
 sky130_fd_sc_hd__or2_1 _23336_ (.A(net159),
    .B(_04779_),
    .X(_04785_));
 sky130_fd_sc_hd__o211a_1 _23337_ (.A1(\top_inst.axis_out_inst.out_buff_data[94] ),
    .A2(_04778_),
    .B1(_04785_),
    .C1(_04782_),
    .X(_01118_));
 sky130_fd_sc_hd__or2_1 _23338_ (.A(net160),
    .B(_04779_),
    .X(_04786_));
 sky130_fd_sc_hd__o211a_1 _23339_ (.A1(net557),
    .A2(_04778_),
    .B1(_04786_),
    .C1(_04782_),
    .X(_01119_));
 sky130_fd_sc_hd__or2_1 _23340_ (.A(net161),
    .B(_04779_),
    .X(_04787_));
 sky130_fd_sc_hd__o211a_1 _23341_ (.A1(net619),
    .A2(_04778_),
    .B1(_04787_),
    .C1(_04782_),
    .X(_01120_));
 sky130_fd_sc_hd__or2_1 _23342_ (.A(net162),
    .B(_04779_),
    .X(_04788_));
 sky130_fd_sc_hd__o211a_1 _23343_ (.A1(net781),
    .A2(_04778_),
    .B1(_04788_),
    .C1(_04782_),
    .X(_01121_));
 sky130_fd_sc_hd__or2_1 _23344_ (.A(net163),
    .B(_04779_),
    .X(_04789_));
 sky130_fd_sc_hd__o211a_1 _23345_ (.A1(net575),
    .A2(_04778_),
    .B1(_04789_),
    .C1(_04782_),
    .X(_01122_));
 sky130_fd_sc_hd__or2_1 _23346_ (.A(net164),
    .B(_04779_),
    .X(_04790_));
 sky130_fd_sc_hd__o211a_1 _23347_ (.A1(net993),
    .A2(_04778_),
    .B1(_04790_),
    .C1(_04782_),
    .X(_01123_));
 sky130_fd_sc_hd__clkbuf_4 _23348_ (.A(_04684_),
    .X(_04791_));
 sky130_fd_sc_hd__buf_2 _23349_ (.A(_04686_),
    .X(_04792_));
 sky130_fd_sc_hd__or2_1 _23350_ (.A(net39),
    .B(_04792_),
    .X(_04793_));
 sky130_fd_sc_hd__o211a_1 _23351_ (.A1(net512),
    .A2(_04791_),
    .B1(_04793_),
    .C1(_04782_),
    .X(_01124_));
 sky130_fd_sc_hd__or2_1 _23352_ (.A(net40),
    .B(_04792_),
    .X(_04794_));
 sky130_fd_sc_hd__clkbuf_4 _23353_ (.A(_04690_),
    .X(_04795_));
 sky130_fd_sc_hd__o211a_1 _23354_ (.A1(net473),
    .A2(_04791_),
    .B1(_04794_),
    .C1(_04795_),
    .X(_01125_));
 sky130_fd_sc_hd__or2_1 _23355_ (.A(net41),
    .B(_04792_),
    .X(_04796_));
 sky130_fd_sc_hd__o211a_1 _23356_ (.A1(net679),
    .A2(_04791_),
    .B1(_04796_),
    .C1(_04795_),
    .X(_01126_));
 sky130_fd_sc_hd__or2_1 _23357_ (.A(net42),
    .B(_04792_),
    .X(_04797_));
 sky130_fd_sc_hd__o211a_1 _23358_ (.A1(net872),
    .A2(_04791_),
    .B1(_04797_),
    .C1(_04795_),
    .X(_01127_));
 sky130_fd_sc_hd__or2_1 _23359_ (.A(net43),
    .B(_04792_),
    .X(_04798_));
 sky130_fd_sc_hd__o211a_1 _23360_ (.A1(net461),
    .A2(_04791_),
    .B1(_04798_),
    .C1(_04795_),
    .X(_01128_));
 sky130_fd_sc_hd__or2_1 _23361_ (.A(net44),
    .B(_04792_),
    .X(_04799_));
 sky130_fd_sc_hd__o211a_1 _23362_ (.A1(net697),
    .A2(_04791_),
    .B1(_04799_),
    .C1(_04795_),
    .X(_01129_));
 sky130_fd_sc_hd__or2_1 _23363_ (.A(net45),
    .B(_04792_),
    .X(_04800_));
 sky130_fd_sc_hd__o211a_1 _23364_ (.A1(net443),
    .A2(_04791_),
    .B1(_04800_),
    .C1(_04795_),
    .X(_01130_));
 sky130_fd_sc_hd__or2_1 _23365_ (.A(net46),
    .B(_04792_),
    .X(_04801_));
 sky130_fd_sc_hd__o211a_1 _23366_ (.A1(net444),
    .A2(_04791_),
    .B1(_04801_),
    .C1(_04795_),
    .X(_01131_));
 sky130_fd_sc_hd__or2_1 _23367_ (.A(net47),
    .B(_04792_),
    .X(_04802_));
 sky130_fd_sc_hd__o211a_1 _23368_ (.A1(net833),
    .A2(_04791_),
    .B1(_04802_),
    .C1(_04795_),
    .X(_01132_));
 sky130_fd_sc_hd__or2_1 _23369_ (.A(net48),
    .B(_04792_),
    .X(_04803_));
 sky130_fd_sc_hd__o211a_1 _23370_ (.A1(net714),
    .A2(_04791_),
    .B1(_04803_),
    .C1(_04795_),
    .X(_01133_));
 sky130_fd_sc_hd__clkbuf_4 _23371_ (.A(_04684_),
    .X(_04804_));
 sky130_fd_sc_hd__buf_2 _23372_ (.A(_04686_),
    .X(_04805_));
 sky130_fd_sc_hd__or2_1 _23373_ (.A(net50),
    .B(_04805_),
    .X(_04806_));
 sky130_fd_sc_hd__o211a_1 _23374_ (.A1(net423),
    .A2(_04804_),
    .B1(_04806_),
    .C1(_04795_),
    .X(_01134_));
 sky130_fd_sc_hd__or2_1 _23375_ (.A(net51),
    .B(_04805_),
    .X(_04807_));
 sky130_fd_sc_hd__clkbuf_4 _23376_ (.A(_04690_),
    .X(_04808_));
 sky130_fd_sc_hd__o211a_1 _23377_ (.A1(net460),
    .A2(_04804_),
    .B1(_04807_),
    .C1(_04808_),
    .X(_01135_));
 sky130_fd_sc_hd__or2_1 _23378_ (.A(net52),
    .B(_04805_),
    .X(_04809_));
 sky130_fd_sc_hd__o211a_1 _23379_ (.A1(net710),
    .A2(_04804_),
    .B1(_04809_),
    .C1(_04808_),
    .X(_01136_));
 sky130_fd_sc_hd__or2_1 _23380_ (.A(net53),
    .B(_04805_),
    .X(_04810_));
 sky130_fd_sc_hd__o211a_1 _23381_ (.A1(net392),
    .A2(_04804_),
    .B1(_04810_),
    .C1(_04808_),
    .X(_01137_));
 sky130_fd_sc_hd__or2_1 _23382_ (.A(net54),
    .B(_04805_),
    .X(_04811_));
 sky130_fd_sc_hd__o211a_1 _23383_ (.A1(net725),
    .A2(_04804_),
    .B1(_04811_),
    .C1(_04808_),
    .X(_01138_));
 sky130_fd_sc_hd__or2_1 _23384_ (.A(net55),
    .B(_04805_),
    .X(_04812_));
 sky130_fd_sc_hd__o211a_1 _23385_ (.A1(net810),
    .A2(_04804_),
    .B1(_04812_),
    .C1(_04808_),
    .X(_01139_));
 sky130_fd_sc_hd__or2_1 _23386_ (.A(net56),
    .B(_04805_),
    .X(_04813_));
 sky130_fd_sc_hd__o211a_1 _23387_ (.A1(net788),
    .A2(_04804_),
    .B1(_04813_),
    .C1(_04808_),
    .X(_01140_));
 sky130_fd_sc_hd__or2_1 _23388_ (.A(net57),
    .B(_04805_),
    .X(_04814_));
 sky130_fd_sc_hd__o211a_1 _23389_ (.A1(net635),
    .A2(_04804_),
    .B1(_04814_),
    .C1(_04808_),
    .X(_01141_));
 sky130_fd_sc_hd__or2_1 _23390_ (.A(net58),
    .B(_04805_),
    .X(_04815_));
 sky130_fd_sc_hd__o211a_1 _23391_ (.A1(net517),
    .A2(_04804_),
    .B1(_04815_),
    .C1(_04808_),
    .X(_01142_));
 sky130_fd_sc_hd__or2_1 _23392_ (.A(net59),
    .B(_04805_),
    .X(_04816_));
 sky130_fd_sc_hd__o211a_1 _23393_ (.A1(net739),
    .A2(_04804_),
    .B1(_04816_),
    .C1(_04808_),
    .X(_01143_));
 sky130_fd_sc_hd__or2_1 _23394_ (.A(net61),
    .B(_04658_),
    .X(_04817_));
 sky130_fd_sc_hd__o211a_1 _23395_ (.A1(net729),
    .A2(_04655_),
    .B1(_04817_),
    .C1(_04808_),
    .X(_01144_));
 sky130_fd_sc_hd__or2_1 _23396_ (.A(net62),
    .B(_04658_),
    .X(_04818_));
 sky130_fd_sc_hd__clkbuf_4 _23397_ (.A(_04869_),
    .X(_04819_));
 sky130_fd_sc_hd__o211a_1 _23398_ (.A1(net842),
    .A2(_04655_),
    .B1(_04818_),
    .C1(_04819_),
    .X(_01145_));
 sky130_fd_sc_hd__or2_1 _23399_ (.A(net63),
    .B(_04658_),
    .X(_04820_));
 sky130_fd_sc_hd__o211a_1 _23400_ (.A1(net451),
    .A2(_04655_),
    .B1(_04820_),
    .C1(_04819_),
    .X(_01146_));
 sky130_fd_sc_hd__or2_1 _23401_ (.A(net64),
    .B(_04658_),
    .X(_04821_));
 sky130_fd_sc_hd__o211a_1 _23402_ (.A1(net410),
    .A2(_04655_),
    .B1(_04821_),
    .C1(_04819_),
    .X(_01147_));
 sky130_fd_sc_hd__or2_1 _23403_ (.A(net65),
    .B(_04658_),
    .X(_04822_));
 sky130_fd_sc_hd__o211a_1 _23404_ (.A1(net801),
    .A2(_04655_),
    .B1(_04822_),
    .C1(_04819_),
    .X(_01148_));
 sky130_fd_sc_hd__or2_1 _23405_ (.A(net66),
    .B(_04658_),
    .X(_04823_));
 sky130_fd_sc_hd__o211a_1 _23406_ (.A1(net751),
    .A2(_04655_),
    .B1(_04823_),
    .C1(_04819_),
    .X(_01149_));
 sky130_fd_sc_hd__or2_1 _23407_ (.A(net67),
    .B(_04658_),
    .X(_04824_));
 sky130_fd_sc_hd__o211a_1 _23408_ (.A1(net623),
    .A2(_04655_),
    .B1(_04824_),
    .C1(_04819_),
    .X(_01150_));
 sky130_fd_sc_hd__or2_1 _23409_ (.A(net68),
    .B(_04658_),
    .X(_04825_));
 sky130_fd_sc_hd__o211a_1 _23410_ (.A1(net530),
    .A2(_04655_),
    .B1(_04825_),
    .C1(_04819_),
    .X(_01151_));
 sky130_fd_sc_hd__o21a_1 _23411_ (.A1(net467),
    .A2(_04856_),
    .B1(_04870_),
    .X(_01152_));
 sky130_fd_sc_hd__or2_1 _23412_ (.A(net619),
    .B(_04596_),
    .X(_04826_));
 sky130_fd_sc_hd__o211a_1 _23413_ (.A1(net1014),
    .A2(_04588_),
    .B1(_04826_),
    .C1(_04819_),
    .X(_01153_));
 sky130_fd_sc_hd__clkbuf_4 _23414_ (.A(_05736_),
    .X(_04827_));
 sky130_fd_sc_hd__or2_1 _23415_ (.A(\top_inst.axis_out_inst.out_buff_data[97] ),
    .B(_04596_),
    .X(_04828_));
 sky130_fd_sc_hd__o211a_1 _23416_ (.A1(net581),
    .A2(_04827_),
    .B1(_04828_),
    .C1(_04819_),
    .X(_01154_));
 sky130_fd_sc_hd__or2_1 _23417_ (.A(\top_inst.axis_out_inst.out_buff_data[98] ),
    .B(_04596_),
    .X(_04829_));
 sky130_fd_sc_hd__o211a_1 _23418_ (.A1(net531),
    .A2(_04827_),
    .B1(_04829_),
    .C1(_04819_),
    .X(_01155_));
 sky130_fd_sc_hd__or2_1 _23419_ (.A(net1107),
    .B(_04596_),
    .X(_04830_));
 sky130_fd_sc_hd__buf_2 _23420_ (.A(_04869_),
    .X(_04831_));
 sky130_fd_sc_hd__o211a_1 _23421_ (.A1(net318),
    .A2(_04827_),
    .B1(_04830_),
    .C1(_04831_),
    .X(_01156_));
 sky130_fd_sc_hd__or2_1 _23422_ (.A(\top_inst.axis_out_inst.out_buff_data[100] ),
    .B(_04596_),
    .X(_04832_));
 sky130_fd_sc_hd__o211a_1 _23423_ (.A1(net371),
    .A2(_04827_),
    .B1(_04832_),
    .C1(_04831_),
    .X(_01157_));
 sky130_fd_sc_hd__or2_1 _23424_ (.A(\top_inst.axis_out_inst.out_buff_data[101] ),
    .B(_04596_),
    .X(_04833_));
 sky130_fd_sc_hd__o211a_1 _23425_ (.A1(net424),
    .A2(_04827_),
    .B1(_04833_),
    .C1(_04831_),
    .X(_01158_));
 sky130_fd_sc_hd__or2_1 _23426_ (.A(\top_inst.axis_out_inst.out_buff_data[102] ),
    .B(_04596_),
    .X(_04834_));
 sky130_fd_sc_hd__o211a_1 _23427_ (.A1(net302),
    .A2(_04827_),
    .B1(_04834_),
    .C1(_04831_),
    .X(_01159_));
 sky130_fd_sc_hd__buf_2 _23428_ (.A(_04863_),
    .X(_04835_));
 sky130_fd_sc_hd__or2_1 _23429_ (.A(\top_inst.axis_out_inst.out_buff_data[103] ),
    .B(_04835_),
    .X(_04836_));
 sky130_fd_sc_hd__o211a_1 _23430_ (.A1(net290),
    .A2(_04827_),
    .B1(_04836_),
    .C1(_04831_),
    .X(_01160_));
 sky130_fd_sc_hd__or2_1 _23431_ (.A(net461),
    .B(_04835_),
    .X(_04837_));
 sky130_fd_sc_hd__o211a_1 _23432_ (.A1(net817),
    .A2(_04827_),
    .B1(_04837_),
    .C1(_04831_),
    .X(_01161_));
 sky130_fd_sc_hd__or2_1 _23433_ (.A(net697),
    .B(_04835_),
    .X(_04838_));
 sky130_fd_sc_hd__o211a_1 _23434_ (.A1(net964),
    .A2(_04827_),
    .B1(_04838_),
    .C1(_04831_),
    .X(_01162_));
 sky130_fd_sc_hd__or2_1 _23435_ (.A(net443),
    .B(_04835_),
    .X(_04839_));
 sky130_fd_sc_hd__o211a_1 _23436_ (.A1(net893),
    .A2(_04827_),
    .B1(_04839_),
    .C1(_04831_),
    .X(_01163_));
 sky130_fd_sc_hd__clkbuf_4 _23437_ (.A(_05736_),
    .X(_04840_));
 sky130_fd_sc_hd__or2_1 _23438_ (.A(net444),
    .B(_04835_),
    .X(_04841_));
 sky130_fd_sc_hd__o211a_1 _23439_ (.A1(net711),
    .A2(_04840_),
    .B1(_04841_),
    .C1(_04831_),
    .X(_01164_));
 sky130_fd_sc_hd__or2_1 _23440_ (.A(\top_inst.axis_out_inst.out_buff_data[108] ),
    .B(_04835_),
    .X(_04842_));
 sky130_fd_sc_hd__o211a_1 _23441_ (.A1(net659),
    .A2(_04840_),
    .B1(_04842_),
    .C1(_04831_),
    .X(_01165_));
 sky130_fd_sc_hd__or2_1 _23442_ (.A(\top_inst.axis_out_inst.out_buff_data[109] ),
    .B(_04835_),
    .X(_04843_));
 sky130_fd_sc_hd__clkbuf_4 _23443_ (.A(_04869_),
    .X(_04844_));
 sky130_fd_sc_hd__o211a_1 _23444_ (.A1(net627),
    .A2(_04840_),
    .B1(_04843_),
    .C1(_04844_),
    .X(_01166_));
 sky130_fd_sc_hd__or2_1 _23445_ (.A(net423),
    .B(_04835_),
    .X(_04845_));
 sky130_fd_sc_hd__o211a_1 _23446_ (.A1(net834),
    .A2(_04840_),
    .B1(_04845_),
    .C1(_04844_),
    .X(_01167_));
 sky130_fd_sc_hd__or2_1 _23447_ (.A(net460),
    .B(_04835_),
    .X(_04846_));
 sky130_fd_sc_hd__o211a_1 _23448_ (.A1(net654),
    .A2(_04840_),
    .B1(_04846_),
    .C1(_04844_),
    .X(_01168_));
 sky130_fd_sc_hd__or2_1 _23449_ (.A(\top_inst.axis_out_inst.out_buff_data[112] ),
    .B(_04835_),
    .X(_04847_));
 sky130_fd_sc_hd__o211a_1 _23450_ (.A1(net508),
    .A2(_04840_),
    .B1(_04847_),
    .C1(_04844_),
    .X(_01169_));
 sky130_fd_sc_hd__or2_1 _23451_ (.A(net392),
    .B(_04864_),
    .X(_04848_));
 sky130_fd_sc_hd__o211a_1 _23452_ (.A1(net923),
    .A2(_04840_),
    .B1(_04848_),
    .C1(_04844_),
    .X(_01170_));
 sky130_fd_sc_hd__or2_1 _23453_ (.A(net725),
    .B(_04864_),
    .X(_04849_));
 sky130_fd_sc_hd__o211a_1 _23454_ (.A1(net740),
    .A2(_04840_),
    .B1(_04849_),
    .C1(_04844_),
    .X(_01171_));
 sky130_fd_sc_hd__or2_1 _23455_ (.A(\top_inst.axis_out_inst.out_buff_data[115] ),
    .B(_04864_),
    .X(_04850_));
 sky130_fd_sc_hd__o211a_1 _23456_ (.A1(net542),
    .A2(_04840_),
    .B1(_04850_),
    .C1(_04844_),
    .X(_01172_));
 sky130_fd_sc_hd__or2_1 _23457_ (.A(\top_inst.axis_out_inst.out_buff_data[116] ),
    .B(_04864_),
    .X(_04851_));
 sky130_fd_sc_hd__o211a_1 _23458_ (.A1(net533),
    .A2(_04840_),
    .B1(_04851_),
    .C1(_04844_),
    .X(_01173_));
 sky130_fd_sc_hd__or2_1 _23459_ (.A(\top_inst.axis_out_inst.out_buff_data[117] ),
    .B(_04864_),
    .X(_04852_));
 sky130_fd_sc_hd__o211a_1 _23460_ (.A1(net260),
    .A2(_04859_),
    .B1(_04852_),
    .C1(_04844_),
    .X(_01174_));
 sky130_fd_sc_hd__or2_1 _23461_ (.A(net517),
    .B(_04864_),
    .X(_04853_));
 sky130_fd_sc_hd__o211a_1 _23462_ (.A1(net884),
    .A2(_04859_),
    .B1(_04853_),
    .C1(_04844_),
    .X(_01175_));
 sky130_fd_sc_hd__or2_1 _23463_ (.A(\top_inst.axis_out_inst.out_buff_data[119] ),
    .B(_04864_),
    .X(_04854_));
 sky130_fd_sc_hd__o211a_1 _23464_ (.A1(net608),
    .A2(_04859_),
    .B1(_04854_),
    .C1(_06180_),
    .X(_01176_));
 sky130_fd_sc_hd__or2_1 _23465_ (.A(\top_inst.axis_out_inst.out_buff_data[120] ),
    .B(_04864_),
    .X(_04855_));
 sky130_fd_sc_hd__o211a_1 _23466_ (.A1(net441),
    .A2(_04859_),
    .B1(_04855_),
    .C1(_06180_),
    .X(_01177_));
 sky130_fd_sc_hd__dfxtp_1 _23467_ (.CLK(clknet_leaf_31_clk),
    .D(net778),
    .Q(\top_inst.axis_out_inst.out_buff_data[121] ));
 sky130_fd_sc_hd__dfxtp_1 _23468_ (.CLK(clknet_leaf_30_clk),
    .D(_00001_),
    .Q(\top_inst.axis_out_inst.out_buff_data[122] ));
 sky130_fd_sc_hd__dfxtp_1 _23469_ (.CLK(clknet_leaf_30_clk),
    .D(_00002_),
    .Q(\top_inst.axis_out_inst.out_buff_data[123] ));
 sky130_fd_sc_hd__dfxtp_1 _23470_ (.CLK(clknet_leaf_32_clk),
    .D(net565),
    .Q(\top_inst.axis_out_inst.out_buff_data[124] ));
 sky130_fd_sc_hd__dfxtp_1 _23471_ (.CLK(clknet_leaf_31_clk),
    .D(net667),
    .Q(\top_inst.axis_out_inst.out_buff_data[125] ));
 sky130_fd_sc_hd__dfxtp_1 _23472_ (.CLK(clknet_leaf_32_clk),
    .D(net472),
    .Q(\top_inst.axis_out_inst.out_buff_data[126] ));
 sky130_fd_sc_hd__dfxtp_1 _23473_ (.CLK(clknet_leaf_30_clk),
    .D(net500),
    .Q(\top_inst.axis_out_inst.out_buff_data[127] ));
 sky130_fd_sc_hd__dfxtp_1 _23474_ (.CLK(clknet_leaf_134_clk),
    .D(net626),
    .Q(\top_inst.axis_out_inst.out_buff_data[64] ));
 sky130_fd_sc_hd__dfxtp_1 _23475_ (.CLK(clknet_leaf_136_clk),
    .D(_00008_),
    .Q(\top_inst.axis_out_inst.out_buff_data[65] ));
 sky130_fd_sc_hd__dfxtp_1 _23476_ (.CLK(clknet_leaf_136_clk),
    .D(_00009_),
    .Q(\top_inst.axis_out_inst.out_buff_data[66] ));
 sky130_fd_sc_hd__dfxtp_1 _23477_ (.CLK(clknet_leaf_136_clk),
    .D(_00010_),
    .Q(\top_inst.axis_out_inst.out_buff_data[67] ));
 sky130_fd_sc_hd__dfxtp_1 _23478_ (.CLK(clknet_leaf_134_clk),
    .D(net349),
    .Q(\top_inst.axis_out_inst.out_buff_data[68] ));
 sky130_fd_sc_hd__dfxtp_1 _23479_ (.CLK(clknet_leaf_134_clk),
    .D(net363),
    .Q(\top_inst.axis_out_inst.out_buff_data[69] ));
 sky130_fd_sc_hd__dfxtp_1 _23480_ (.CLK(clknet_leaf_136_clk),
    .D(net361),
    .Q(\top_inst.axis_out_inst.out_buff_data[70] ));
 sky130_fd_sc_hd__dfxtp_1 _23481_ (.CLK(clknet_leaf_136_clk),
    .D(net338),
    .Q(\top_inst.axis_out_inst.out_buff_data[71] ));
 sky130_fd_sc_hd__dfxtp_1 _23482_ (.CLK(clknet_leaf_137_clk),
    .D(_00015_),
    .Q(\top_inst.axis_out_inst.out_buff_data[72] ));
 sky130_fd_sc_hd__dfxtp_1 _23483_ (.CLK(clknet_leaf_134_clk),
    .D(net368),
    .Q(\top_inst.axis_out_inst.out_buff_data[73] ));
 sky130_fd_sc_hd__dfxtp_1 _23484_ (.CLK(clknet_leaf_137_clk),
    .D(_00017_),
    .Q(\top_inst.axis_out_inst.out_buff_data[74] ));
 sky130_fd_sc_hd__dfxtp_1 _23485_ (.CLK(clknet_leaf_138_clk),
    .D(_00018_),
    .Q(\top_inst.axis_out_inst.out_buff_data[75] ));
 sky130_fd_sc_hd__dfxtp_1 _23486_ (.CLK(clknet_leaf_138_clk),
    .D(_00019_),
    .Q(\top_inst.axis_out_inst.out_buff_data[76] ));
 sky130_fd_sc_hd__dfxtp_1 _23487_ (.CLK(clknet_leaf_141_clk),
    .D(_00020_),
    .Q(\top_inst.axis_out_inst.out_buff_data[77] ));
 sky130_fd_sc_hd__dfxtp_1 _23488_ (.CLK(clknet_leaf_140_clk),
    .D(net571),
    .Q(\top_inst.axis_out_inst.out_buff_data[78] ));
 sky130_fd_sc_hd__dfxtp_1 _23489_ (.CLK(clknet_leaf_140_clk),
    .D(net615),
    .Q(\top_inst.axis_out_inst.out_buff_data[79] ));
 sky130_fd_sc_hd__dfxtp_1 _23490_ (.CLK(clknet_leaf_140_clk),
    .D(net641),
    .Q(\top_inst.axis_out_inst.out_buff_data[80] ));
 sky130_fd_sc_hd__dfxtp_1 _23491_ (.CLK(clknet_leaf_139_clk),
    .D(_00024_),
    .Q(\top_inst.axis_out_inst.out_buff_data[81] ));
 sky130_fd_sc_hd__dfxtp_1 _23492_ (.CLK(clknet_leaf_140_clk),
    .D(net523),
    .Q(\top_inst.axis_out_inst.out_buff_data[82] ));
 sky130_fd_sc_hd__dfxtp_1 _23493_ (.CLK(clknet_leaf_142_clk),
    .D(_00026_),
    .Q(\top_inst.axis_out_inst.out_buff_data[83] ));
 sky130_fd_sc_hd__dfxtp_1 _23494_ (.CLK(clknet_leaf_143_clk),
    .D(_00027_),
    .Q(\top_inst.axis_out_inst.out_buff_data[84] ));
 sky130_fd_sc_hd__dfxtp_1 _23495_ (.CLK(clknet_leaf_143_clk),
    .D(_00028_),
    .Q(\top_inst.axis_out_inst.out_buff_data[85] ));
 sky130_fd_sc_hd__dfxtp_1 _23496_ (.CLK(clknet_leaf_140_clk),
    .D(net475),
    .Q(\top_inst.axis_out_inst.out_buff_data[86] ));
 sky130_fd_sc_hd__dfxtp_1 _23497_ (.CLK(clknet_leaf_142_clk),
    .D(_00030_),
    .Q(\top_inst.axis_out_inst.out_buff_data[87] ));
 sky130_fd_sc_hd__dfxtp_1 _23498_ (.CLK(clknet_leaf_140_clk),
    .D(_00031_),
    .Q(\top_inst.axis_out_inst.out_buff_data[88] ));
 sky130_fd_sc_hd__dfxtp_1 _23499_ (.CLK(clknet_leaf_141_clk),
    .D(_00032_),
    .Q(\top_inst.axis_out_inst.out_buff_data[89] ));
 sky130_fd_sc_hd__dfxtp_1 _23500_ (.CLK(clknet_leaf_139_clk),
    .D(_00033_),
    .Q(\top_inst.axis_out_inst.out_buff_data[90] ));
 sky130_fd_sc_hd__dfxtp_1 _23501_ (.CLK(clknet_leaf_140_clk),
    .D(_00034_),
    .Q(\top_inst.axis_out_inst.out_buff_data[91] ));
 sky130_fd_sc_hd__dfxtp_1 _23502_ (.CLK(clknet_leaf_141_clk),
    .D(_00035_),
    .Q(\top_inst.axis_out_inst.out_buff_data[92] ));
 sky130_fd_sc_hd__dfxtp_1 _23503_ (.CLK(clknet_leaf_140_clk),
    .D(net685),
    .Q(\top_inst.axis_out_inst.out_buff_data[93] ));
 sky130_fd_sc_hd__dfxtp_2 _23504_ (.CLK(clknet_leaf_139_clk),
    .D(_00037_),
    .Q(\top_inst.axis_out_inst.out_buff_data[94] ));
 sky130_fd_sc_hd__dfxtp_1 _23505_ (.CLK(clknet_leaf_134_clk),
    .D(net429),
    .Q(\top_inst.axis_out_inst.out_buff_data[95] ));
 sky130_fd_sc_hd__dfxtp_1 _23506_ (.CLK(clknet_leaf_134_clk),
    .D(net455),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _23507_ (.CLK(clknet_leaf_136_clk),
    .D(net326),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _23508_ (.CLK(clknet_leaf_135_clk),
    .D(net283),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _23509_ (.CLK(clknet_leaf_136_clk),
    .D(net314),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _23510_ (.CLK(clknet_leaf_137_clk),
    .D(_00043_),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _23511_ (.CLK(clknet_leaf_137_clk),
    .D(_00044_),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _23512_ (.CLK(clknet_leaf_137_clk),
    .D(_00045_),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _23513_ (.CLK(clknet_leaf_137_clk),
    .D(_00046_),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _23514_ (.CLK(clknet_leaf_137_clk),
    .D(_00047_),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _23515_ (.CLK(clknet_leaf_137_clk),
    .D(_00048_),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _23516_ (.CLK(clknet_leaf_138_clk),
    .D(_00049_),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _23517_ (.CLK(clknet_leaf_138_clk),
    .D(net754),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _23518_ (.CLK(clknet_leaf_138_clk),
    .D(net840),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _23519_ (.CLK(clknet_leaf_138_clk),
    .D(net819),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _23520_ (.CLK(clknet_leaf_138_clk),
    .D(_00053_),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _23521_ (.CLK(clknet_leaf_139_clk),
    .D(net545),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _23522_ (.CLK(clknet_leaf_139_clk),
    .D(net412),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _23523_ (.CLK(clknet_leaf_138_clk),
    .D(_00056_),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _23524_ (.CLK(clknet_leaf_139_clk),
    .D(net504),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _23525_ (.CLK(clknet_leaf_1_clk),
    .D(_00058_),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _23526_ (.CLK(clknet_leaf_1_clk),
    .D(net887),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _23527_ (.CLK(clknet_leaf_139_clk),
    .D(net649),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _23528_ (.CLK(clknet_leaf_139_clk),
    .D(_00061_),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _23529_ (.CLK(clknet_leaf_139_clk),
    .D(net671),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _23530_ (.CLK(clknet_leaf_140_clk),
    .D(net525),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _23531_ (.CLK(clknet_leaf_142_clk),
    .D(_00064_),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _23532_ (.CLK(clknet_leaf_139_clk),
    .D(net431),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _23533_ (.CLK(clknet_leaf_140_clk),
    .D(net683),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _23534_ (.CLK(clknet_leaf_140_clk),
    .D(net669),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _23535_ (.CLK(clknet_leaf_140_clk),
    .D(net562),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _23536_ (.CLK(clknet_leaf_139_clk),
    .D(_00069_),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _23537_ (.CLK(clknet_leaf_141_clk),
    .D(_00070_),
    .Q(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _23538_ (.CLK(clknet_leaf_132_clk),
    .D(_00071_),
    .Q(\top_inst.axis_out_inst.out_buff_data[32] ));
 sky130_fd_sc_hd__dfxtp_1 _23539_ (.CLK(clknet_leaf_131_clk),
    .D(_00072_),
    .Q(\top_inst.axis_out_inst.out_buff_data[33] ));
 sky130_fd_sc_hd__dfxtp_1 _23540_ (.CLK(clknet_leaf_128_clk),
    .D(net482),
    .Q(\top_inst.axis_out_inst.out_buff_data[34] ));
 sky130_fd_sc_hd__dfxtp_1 _23541_ (.CLK(clknet_leaf_128_clk),
    .D(net479),
    .Q(\top_inst.axis_out_inst.out_buff_data[35] ));
 sky130_fd_sc_hd__dfxtp_1 _23542_ (.CLK(clknet_leaf_129_clk),
    .D(_00075_),
    .Q(\top_inst.axis_out_inst.out_buff_data[36] ));
 sky130_fd_sc_hd__dfxtp_1 _23543_ (.CLK(clknet_leaf_130_clk),
    .D(_00076_),
    .Q(\top_inst.axis_out_inst.out_buff_data[37] ));
 sky130_fd_sc_hd__dfxtp_1 _23544_ (.CLK(clknet_leaf_130_clk),
    .D(_00077_),
    .Q(\top_inst.axis_out_inst.out_buff_data[38] ));
 sky130_fd_sc_hd__dfxtp_1 _23545_ (.CLK(clknet_leaf_129_clk),
    .D(_00078_),
    .Q(\top_inst.axis_out_inst.out_buff_data[39] ));
 sky130_fd_sc_hd__dfxtp_1 _23546_ (.CLK(clknet_leaf_129_clk),
    .D(_00079_),
    .Q(\top_inst.axis_out_inst.out_buff_data[40] ));
 sky130_fd_sc_hd__dfxtp_1 _23547_ (.CLK(clknet_leaf_103_clk),
    .D(net521),
    .Q(\top_inst.axis_out_inst.out_buff_data[41] ));
 sky130_fd_sc_hd__dfxtp_1 _23548_ (.CLK(clknet_leaf_130_clk),
    .D(_00081_),
    .Q(\top_inst.axis_out_inst.out_buff_data[42] ));
 sky130_fd_sc_hd__dfxtp_1 _23549_ (.CLK(clknet_leaf_131_clk),
    .D(_00082_),
    .Q(\top_inst.axis_out_inst.out_buff_data[43] ));
 sky130_fd_sc_hd__dfxtp_1 _23550_ (.CLK(clknet_leaf_130_clk),
    .D(_00083_),
    .Q(\top_inst.axis_out_inst.out_buff_data[44] ));
 sky130_fd_sc_hd__dfxtp_1 _23551_ (.CLK(clknet_leaf_102_clk),
    .D(net550),
    .Q(\top_inst.axis_out_inst.out_buff_data[45] ));
 sky130_fd_sc_hd__dfxtp_1 _23552_ (.CLK(clknet_leaf_129_clk),
    .D(_00085_),
    .Q(\top_inst.axis_out_inst.out_buff_data[46] ));
 sky130_fd_sc_hd__dfxtp_1 _23553_ (.CLK(clknet_leaf_105_clk),
    .D(_00086_),
    .Q(\top_inst.axis_out_inst.out_buff_data[47] ));
 sky130_fd_sc_hd__dfxtp_1 _23554_ (.CLK(clknet_leaf_129_clk),
    .D(_00087_),
    .Q(\top_inst.axis_out_inst.out_buff_data[48] ));
 sky130_fd_sc_hd__dfxtp_1 _23555_ (.CLK(clknet_leaf_102_clk),
    .D(_00088_),
    .Q(\top_inst.axis_out_inst.out_buff_data[49] ));
 sky130_fd_sc_hd__dfxtp_1 _23556_ (.CLK(clknet_leaf_102_clk),
    .D(_00089_),
    .Q(\top_inst.axis_out_inst.out_buff_data[50] ));
 sky130_fd_sc_hd__dfxtp_1 _23557_ (.CLK(clknet_leaf_102_clk),
    .D(_00090_),
    .Q(\top_inst.axis_out_inst.out_buff_data[51] ));
 sky130_fd_sc_hd__dfxtp_1 _23558_ (.CLK(clknet_leaf_102_clk),
    .D(net915),
    .Q(\top_inst.axis_out_inst.out_buff_data[52] ));
 sky130_fd_sc_hd__dfxtp_1 _23559_ (.CLK(clknet_leaf_100_clk),
    .D(net806),
    .Q(\top_inst.axis_out_inst.out_buff_data[53] ));
 sky130_fd_sc_hd__dfxtp_1 _23560_ (.CLK(clknet_leaf_100_clk),
    .D(_00093_),
    .Q(\top_inst.axis_out_inst.out_buff_data[54] ));
 sky130_fd_sc_hd__dfxtp_1 _23561_ (.CLK(clknet_leaf_103_clk),
    .D(net701),
    .Q(\top_inst.axis_out_inst.out_buff_data[55] ));
 sky130_fd_sc_hd__dfxtp_1 _23562_ (.CLK(clknet_leaf_100_clk),
    .D(net815),
    .Q(\top_inst.axis_out_inst.out_buff_data[56] ));
 sky130_fd_sc_hd__dfxtp_1 _23563_ (.CLK(clknet_leaf_100_clk),
    .D(net792),
    .Q(\top_inst.axis_out_inst.out_buff_data[57] ));
 sky130_fd_sc_hd__dfxtp_1 _23564_ (.CLK(clknet_leaf_102_clk),
    .D(_00097_),
    .Q(\top_inst.axis_out_inst.out_buff_data[58] ));
 sky130_fd_sc_hd__dfxtp_1 _23565_ (.CLK(clknet_leaf_100_clk),
    .D(net721),
    .Q(\top_inst.axis_out_inst.out_buff_data[59] ));
 sky130_fd_sc_hd__dfxtp_1 _23566_ (.CLK(clknet_leaf_103_clk),
    .D(net552),
    .Q(\top_inst.axis_out_inst.out_buff_data[60] ));
 sky130_fd_sc_hd__dfxtp_1 _23567_ (.CLK(clknet_leaf_103_clk),
    .D(_00100_),
    .Q(\top_inst.axis_out_inst.out_buff_data[61] ));
 sky130_fd_sc_hd__dfxtp_1 _23568_ (.CLK(clknet_leaf_103_clk),
    .D(_00101_),
    .Q(\top_inst.axis_out_inst.out_buff_data[62] ));
 sky130_fd_sc_hd__dfxtp_1 _23569_ (.CLK(clknet_leaf_103_clk),
    .D(_00102_),
    .Q(\top_inst.axis_out_inst.out_buff_data[63] ));
 sky130_fd_sc_hd__dfxtp_1 _23570_ (.CLK(clknet_leaf_104_clk),
    .D(net738),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _23571_ (.CLK(clknet_leaf_107_clk),
    .D(_00104_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _23572_ (.CLK(clknet_leaf_108_clk),
    .D(_00105_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _23573_ (.CLK(clknet_leaf_129_clk),
    .D(_00106_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _23574_ (.CLK(clknet_leaf_108_clk),
    .D(net498),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _23575_ (.CLK(clknet_leaf_104_clk),
    .D(_00108_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _23576_ (.CLK(clknet_leaf_107_clk),
    .D(_00109_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _23577_ (.CLK(clknet_leaf_107_clk),
    .D(_00110_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _23578_ (.CLK(clknet_leaf_107_clk),
    .D(_00111_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _23579_ (.CLK(clknet_leaf_106_clk),
    .D(_00112_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _23580_ (.CLK(clknet_leaf_106_clk),
    .D(_00113_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _23581_ (.CLK(clknet_leaf_107_clk),
    .D(_00114_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _23582_ (.CLK(clknet_leaf_106_clk),
    .D(_00115_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _23583_ (.CLK(clknet_leaf_110_clk),
    .D(_00116_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _23584_ (.CLK(clknet_leaf_106_clk),
    .D(net316),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _23585_ (.CLK(clknet_leaf_106_clk),
    .D(net279),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _23586_ (.CLK(clknet_leaf_106_clk),
    .D(net271),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _23587_ (.CLK(clknet_leaf_105_clk),
    .D(net281),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _23588_ (.CLK(clknet_leaf_106_clk),
    .D(net269),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _23589_ (.CLK(clknet_4_8__leaf_clk),
    .D(_00122_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _23590_ (.CLK(clknet_leaf_101_clk),
    .D(_00123_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _23591_ (.CLK(clknet_leaf_101_clk),
    .D(_00124_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _23592_ (.CLK(clknet_leaf_101_clk),
    .D(_00125_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _23593_ (.CLK(clknet_leaf_101_clk),
    .D(_00126_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _23594_ (.CLK(clknet_leaf_101_clk),
    .D(_00127_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _23595_ (.CLK(clknet_leaf_100_clk),
    .D(_00128_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _23596_ (.CLK(clknet_leaf_100_clk),
    .D(_00129_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _23597_ (.CLK(clknet_leaf_101_clk),
    .D(_00130_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _23598_ (.CLK(clknet_leaf_101_clk),
    .D(_00131_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _23599_ (.CLK(clknet_leaf_103_clk),
    .D(net328),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _23600_ (.CLK(clknet_leaf_103_clk),
    .D(net560),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _23601_ (.CLK(clknet_leaf_103_clk),
    .D(net519),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _23602_ (.CLK(clknet_leaf_104_clk),
    .D(_00135_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _23603_ (.CLK(clknet_leaf_103_clk),
    .D(net448),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _23604_ (.CLK(clknet_leaf_104_clk),
    .D(_00137_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _23605_ (.CLK(clknet_leaf_104_clk),
    .D(_00138_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _23606_ (.CLK(clknet_leaf_104_clk),
    .D(_00139_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _23607_ (.CLK(clknet_leaf_104_clk),
    .D(net798),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _23608_ (.CLK(clknet_leaf_103_clk),
    .D(net459),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _23609_ (.CLK(clknet_leaf_104_clk),
    .D(net547),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _23610_ (.CLK(clknet_leaf_104_clk),
    .D(net446),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _23611_ (.CLK(clknet_leaf_104_clk),
    .D(_00144_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _23612_ (.CLK(clknet_leaf_105_clk),
    .D(_00145_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _23613_ (.CLK(clknet_leaf_105_clk),
    .D(_00146_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _23614_ (.CLK(clknet_leaf_105_clk),
    .D(_00147_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _23615_ (.CLK(clknet_leaf_105_clk),
    .D(net273),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _23616_ (.CLK(clknet_leaf_105_clk),
    .D(net539),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _23617_ (.CLK(clknet_leaf_105_clk),
    .D(net588),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _23618_ (.CLK(clknet_leaf_105_clk),
    .D(net574),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _23619_ (.CLK(clknet_leaf_102_clk),
    .D(net502),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _23620_ (.CLK(clknet_leaf_102_clk),
    .D(net487),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _23621_ (.CLK(clknet_leaf_102_clk),
    .D(net255),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _23622_ (.CLK(clknet_leaf_102_clk),
    .D(net263),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _23623_ (.CLK(clknet_leaf_100_clk),
    .D(net470),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _23624_ (.CLK(clknet_leaf_100_clk),
    .D(net511),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _23625_ (.CLK(clknet_leaf_102_clk),
    .D(net265),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _23626_ (.CLK(clknet_leaf_100_clk),
    .D(net386),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _23627_ (.CLK(clknet_leaf_100_clk),
    .D(_00160_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _23628_ (.CLK(clknet_leaf_102_clk),
    .D(net275),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _23629_ (.CLK(clknet_leaf_102_clk),
    .D(net257),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _23630_ (.CLK(clknet_leaf_102_clk),
    .D(net267),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _23631_ (.CLK(clknet_leaf_102_clk),
    .D(net507),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _23632_ (.CLK(clknet_leaf_103_clk),
    .D(_00165_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _23633_ (.CLK(clknet_leaf_103_clk),
    .D(_00166_),
    .Q(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _23634_ (.CLK(clknet_leaf_125_clk),
    .D(net931),
    .Q(\top_inst.axis_out_inst.out_buff_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _23635_ (.CLK(clknet_leaf_108_clk),
    .D(net433),
    .Q(\top_inst.axis_out_inst.out_buff_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _23636_ (.CLK(clknet_leaf_125_clk),
    .D(_00169_),
    .Q(\top_inst.axis_out_inst.out_buff_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _23637_ (.CLK(clknet_leaf_126_clk),
    .D(_00170_),
    .Q(\top_inst.axis_out_inst.out_buff_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _23638_ (.CLK(clknet_leaf_108_clk),
    .D(net399),
    .Q(\top_inst.axis_out_inst.out_buff_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _23639_ (.CLK(clknet_leaf_126_clk),
    .D(_00172_),
    .Q(\top_inst.axis_out_inst.out_buff_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23640_ (.CLK(clknet_leaf_126_clk),
    .D(net403),
    .Q(\top_inst.axis_out_inst.out_buff_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _23641_ (.CLK(clknet_leaf_125_clk),
    .D(net419),
    .Q(\top_inst.axis_out_inst.out_buff_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _23642_ (.CLK(clknet_leaf_127_clk),
    .D(_00175_),
    .Q(\top_inst.axis_out_inst.out_buff_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _23643_ (.CLK(clknet_leaf_126_clk),
    .D(net374),
    .Q(\top_inst.axis_out_inst.out_buff_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _23644_ (.CLK(clknet_leaf_126_clk),
    .D(net358),
    .Q(\top_inst.axis_out_inst.out_buff_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _23645_ (.CLK(clknet_leaf_123_clk),
    .D(net593),
    .Q(\top_inst.axis_out_inst.out_buff_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _23646_ (.CLK(clknet_leaf_127_clk),
    .D(_00179_),
    .Q(\top_inst.axis_out_inst.out_buff_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _23647_ (.CLK(clknet_leaf_127_clk),
    .D(_00180_),
    .Q(\top_inst.axis_out_inst.out_buff_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _23648_ (.CLK(clknet_leaf_127_clk),
    .D(_00181_),
    .Q(\top_inst.axis_out_inst.out_buff_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _23649_ (.CLK(clknet_leaf_128_clk),
    .D(net324),
    .Q(\top_inst.axis_out_inst.out_buff_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _23650_ (.CLK(clknet_leaf_132_clk),
    .D(net347),
    .Q(\top_inst.axis_out_inst.out_buff_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _23651_ (.CLK(clknet_leaf_122_clk),
    .D(_00184_),
    .Q(\top_inst.axis_out_inst.out_buff_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _23652_ (.CLK(clknet_leaf_128_clk),
    .D(net342),
    .Q(\top_inst.axis_out_inst.out_buff_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _23653_ (.CLK(clknet_leaf_128_clk),
    .D(net351),
    .Q(\top_inst.axis_out_inst.out_buff_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _23654_ (.CLK(clknet_leaf_135_clk),
    .D(_00187_),
    .Q(\top_inst.axis_out_inst.out_buff_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _23655_ (.CLK(clknet_leaf_135_clk),
    .D(_00188_),
    .Q(\top_inst.axis_out_inst.out_buff_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _23656_ (.CLK(clknet_leaf_132_clk),
    .D(net353),
    .Q(\top_inst.axis_out_inst.out_buff_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _23657_ (.CLK(clknet_leaf_132_clk),
    .D(net366),
    .Q(\top_inst.axis_out_inst.out_buff_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _23658_ (.CLK(clknet_leaf_135_clk),
    .D(_00191_),
    .Q(\top_inst.axis_out_inst.out_buff_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _23659_ (.CLK(clknet_leaf_132_clk),
    .D(net527),
    .Q(\top_inst.axis_out_inst.out_buff_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _23660_ (.CLK(clknet_leaf_135_clk),
    .D(_00193_),
    .Q(\top_inst.axis_out_inst.out_buff_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _23661_ (.CLK(clknet_leaf_135_clk),
    .D(_00194_),
    .Q(\top_inst.axis_out_inst.out_buff_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _23662_ (.CLK(clknet_leaf_132_clk),
    .D(net309),
    .Q(\top_inst.axis_out_inst.out_buff_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _23663_ (.CLK(clknet_leaf_132_clk),
    .D(net376),
    .Q(\top_inst.axis_out_inst.out_buff_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _23664_ (.CLK(clknet_leaf_132_clk),
    .D(net340),
    .Q(\top_inst.axis_out_inst.out_buff_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _23665_ (.CLK(clknet_leaf_132_clk),
    .D(net384),
    .Q(\top_inst.axis_out_inst.out_buff_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _23666_ (.CLK(clknet_leaf_124_clk),
    .D(_00199_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _23667_ (.CLK(clknet_leaf_124_clk),
    .D(_00200_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _23668_ (.CLK(clknet_leaf_125_clk),
    .D(net409),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _23669_ (.CLK(clknet_leaf_116_clk),
    .D(net344),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _23670_ (.CLK(clknet_leaf_116_clk),
    .D(net356),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _23671_ (.CLK(clknet_leaf_116_clk),
    .D(net813),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _23672_ (.CLK(clknet_leaf_116_clk),
    .D(_00205_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _23673_ (.CLK(clknet_leaf_116_clk),
    .D(_00206_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _23674_ (.CLK(clknet_leaf_116_clk),
    .D(net847),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _23675_ (.CLK(clknet_leaf_116_clk),
    .D(net465),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _23676_ (.CLK(clknet_leaf_116_clk),
    .D(net427),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _23677_ (.CLK(clknet_leaf_116_clk),
    .D(net421),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _23678_ (.CLK(clknet_leaf_117_clk),
    .D(net827),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _23679_ (.CLK(clknet_leaf_116_clk),
    .D(net597),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _23680_ (.CLK(clknet_leaf_117_clk),
    .D(net484),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _23681_ (.CLK(clknet_leaf_117_clk),
    .D(net438),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _23682_ (.CLK(clknet_leaf_117_clk),
    .D(net312),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _23683_ (.CLK(clknet_leaf_119_clk),
    .D(_00216_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _23684_ (.CLK(clknet_leaf_117_clk),
    .D(net436),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _23685_ (.CLK(clknet_leaf_118_clk),
    .D(_00218_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _23686_ (.CLK(clknet_leaf_118_clk),
    .D(_00219_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _23687_ (.CLK(clknet_leaf_119_clk),
    .D(_00220_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _23688_ (.CLK(clknet_leaf_119_clk),
    .D(_00221_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _23689_ (.CLK(clknet_leaf_119_clk),
    .D(_00222_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _23690_ (.CLK(clknet_leaf_120_clk),
    .D(_00223_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _23691_ (.CLK(clknet_leaf_120_clk),
    .D(_00224_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _23692_ (.CLK(clknet_leaf_120_clk),
    .D(_00225_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _23693_ (.CLK(clknet_leaf_119_clk),
    .D(_00226_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _23694_ (.CLK(clknet_leaf_119_clk),
    .D(_00227_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _23695_ (.CLK(clknet_leaf_119_clk),
    .D(_00228_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _23696_ (.CLK(clknet_leaf_120_clk),
    .D(net401),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _23697_ (.CLK(clknet_leaf_121_clk),
    .D(net491),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _23698_ (.CLK(clknet_leaf_124_clk),
    .D(_00231_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _23699_ (.CLK(clknet_leaf_124_clk),
    .D(_00232_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _23700_ (.CLK(clknet_leaf_125_clk),
    .D(_00233_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _23701_ (.CLK(clknet_leaf_125_clk),
    .D(_00234_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _23702_ (.CLK(clknet_leaf_125_clk),
    .D(net601),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _23703_ (.CLK(clknet_leaf_116_clk),
    .D(_00236_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _23704_ (.CLK(clknet_leaf_125_clk),
    .D(net555),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _23705_ (.CLK(clknet_leaf_125_clk),
    .D(net529),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _23706_ (.CLK(clknet_leaf_124_clk),
    .D(_00239_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _23707_ (.CLK(clknet_leaf_124_clk),
    .D(_00240_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _23708_ (.CLK(clknet_leaf_124_clk),
    .D(_00241_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _23709_ (.CLK(clknet_leaf_124_clk),
    .D(_00242_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _23710_ (.CLK(clknet_leaf_123_clk),
    .D(_00243_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _23711_ (.CLK(clknet_leaf_124_clk),
    .D(_00244_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _23712_ (.CLK(clknet_leaf_123_clk),
    .D(_00245_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _23713_ (.CLK(clknet_leaf_123_clk),
    .D(_00246_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _23714_ (.CLK(clknet_leaf_123_clk),
    .D(_00247_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _23715_ (.CLK(clknet_leaf_121_clk),
    .D(_00248_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _23716_ (.CLK(clknet_leaf_121_clk),
    .D(_00249_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _23717_ (.CLK(clknet_leaf_121_clk),
    .D(_00250_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _23718_ (.CLK(clknet_leaf_120_clk),
    .D(_00251_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _23719_ (.CLK(clknet_leaf_120_clk),
    .D(_00252_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _23720_ (.CLK(clknet_leaf_121_clk),
    .D(_00253_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _23721_ (.CLK(clknet_leaf_121_clk),
    .D(_00254_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _23722_ (.CLK(clknet_leaf_120_clk),
    .D(_00255_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _23723_ (.CLK(clknet_leaf_120_clk),
    .D(_00256_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _23724_ (.CLK(clknet_leaf_120_clk),
    .D(_00257_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _23725_ (.CLK(clknet_leaf_136_clk),
    .D(net307),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _23726_ (.CLK(clknet_leaf_121_clk),
    .D(_00259_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _23727_ (.CLK(clknet_leaf_121_clk),
    .D(_00260_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _23728_ (.CLK(clknet_leaf_121_clk),
    .D(_00261_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _23729_ (.CLK(clknet_leaf_121_clk),
    .D(_00262_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _23730_ (.CLK(clknet_leaf_125_clk),
    .D(net496),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _23731_ (.CLK(clknet_leaf_125_clk),
    .D(_00264_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _23732_ (.CLK(clknet_leaf_125_clk),
    .D(_00265_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _23733_ (.CLK(clknet_leaf_126_clk),
    .D(net457),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _23734_ (.CLK(clknet_leaf_125_clk),
    .D(_00267_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _23735_ (.CLK(clknet_leaf_126_clk),
    .D(net453),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _23736_ (.CLK(clknet_leaf_125_clk),
    .D(_00269_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _23737_ (.CLK(clknet_leaf_127_clk),
    .D(_00270_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _23738_ (.CLK(clknet_leaf_127_clk),
    .D(net569),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _23739_ (.CLK(clknet_leaf_127_clk),
    .D(_00272_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _23740_ (.CLK(clknet_leaf_127_clk),
    .D(_00273_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _23741_ (.CLK(clknet_leaf_122_clk),
    .D(net536),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _23742_ (.CLK(clknet_leaf_127_clk),
    .D(net450),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _23743_ (.CLK(clknet_leaf_122_clk),
    .D(_00276_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _23744_ (.CLK(clknet_leaf_127_clk),
    .D(net516),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _23745_ (.CLK(clknet_leaf_122_clk),
    .D(_00278_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _23746_ (.CLK(clknet_leaf_122_clk),
    .D(_00279_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _23747_ (.CLK(clknet_leaf_122_clk),
    .D(net320),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _23748_ (.CLK(clknet_leaf_122_clk),
    .D(_00281_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _23749_ (.CLK(clknet_leaf_122_clk),
    .D(net330),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _23750_ (.CLK(clknet_leaf_135_clk),
    .D(net293),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _23751_ (.CLK(clknet_leaf_135_clk),
    .D(net299),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _23752_ (.CLK(clknet_leaf_122_clk),
    .D(net334),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _23753_ (.CLK(clknet_leaf_122_clk),
    .D(net322),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _23754_ (.CLK(clknet_leaf_135_clk),
    .D(net287),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _23755_ (.CLK(clknet_leaf_135_clk),
    .D(net277),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _23756_ (.CLK(clknet_leaf_135_clk),
    .D(net289),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _23757_ (.CLK(clknet_leaf_135_clk),
    .D(net370),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _23758_ (.CLK(clknet_leaf_121_clk),
    .D(_00291_),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _23759_ (.CLK(clknet_leaf_122_clk),
    .D(net305),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _23760_ (.CLK(clknet_leaf_123_clk),
    .D(net336),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _23761_ (.CLK(clknet_leaf_122_clk),
    .D(net301),
    .Q(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][31] ));
 sky130_fd_sc_hd__dfxtp_2 _23762_ (.CLK(clknet_leaf_66_clk),
    .D(_00295_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _23763_ (.CLK(clknet_leaf_66_clk),
    .D(_00296_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _23764_ (.CLK(clknet_leaf_66_clk),
    .D(_00297_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _23765_ (.CLK(clknet_leaf_66_clk),
    .D(_00298_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _23766_ (.CLK(clknet_leaf_66_clk),
    .D(_00299_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _23767_ (.CLK(clknet_leaf_66_clk),
    .D(_00300_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23768_ (.CLK(clknet_leaf_66_clk),
    .D(_00301_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _23769_ (.CLK(clknet_leaf_66_clk),
    .D(_00302_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _23770_ (.CLK(clknet_leaf_62_clk),
    .D(_00303_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[0] ));
 sky130_fd_sc_hd__dfxtp_1 _23771_ (.CLK(clknet_leaf_62_clk),
    .D(_00304_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[1] ));
 sky130_fd_sc_hd__dfxtp_1 _23772_ (.CLK(clknet_leaf_63_clk),
    .D(_00305_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _23773_ (.CLK(clknet_leaf_63_clk),
    .D(_00306_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[3] ));
 sky130_fd_sc_hd__dfxtp_1 _23774_ (.CLK(clknet_leaf_63_clk),
    .D(_00307_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[4] ));
 sky130_fd_sc_hd__dfxtp_1 _23775_ (.CLK(clknet_leaf_63_clk),
    .D(_00308_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23776_ (.CLK(clknet_leaf_64_clk),
    .D(_00309_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[6] ));
 sky130_fd_sc_hd__dfxtp_1 _23777_ (.CLK(clknet_leaf_64_clk),
    .D(_00310_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[7] ));
 sky130_fd_sc_hd__dfxtp_1 _23778_ (.CLK(clknet_leaf_64_clk),
    .D(_00311_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[8] ));
 sky130_fd_sc_hd__dfxtp_1 _23779_ (.CLK(clknet_leaf_65_clk),
    .D(_00312_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[9] ));
 sky130_fd_sc_hd__dfxtp_1 _23780_ (.CLK(clknet_leaf_65_clk),
    .D(_00313_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[10] ));
 sky130_fd_sc_hd__dfxtp_1 _23781_ (.CLK(clknet_leaf_65_clk),
    .D(_00314_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[11] ));
 sky130_fd_sc_hd__dfxtp_1 _23782_ (.CLK(clknet_leaf_65_clk),
    .D(_00315_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[12] ));
 sky130_fd_sc_hd__dfxtp_1 _23783_ (.CLK(clknet_leaf_65_clk),
    .D(_00316_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _23784_ (.CLK(clknet_leaf_65_clk),
    .D(_00317_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[14] ));
 sky130_fd_sc_hd__dfxtp_1 _23785_ (.CLK(clknet_leaf_65_clk),
    .D(_00318_),
    .Q(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[15] ));
 sky130_fd_sc_hd__dfxtp_1 _23786_ (.CLK(clknet_leaf_70_clk),
    .D(_00319_),
    .Q(\top_inst.grid_inst.data_path_wires[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _23787_ (.CLK(clknet_leaf_70_clk),
    .D(_00320_),
    .Q(\top_inst.grid_inst.data_path_wires[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _23788_ (.CLK(clknet_leaf_70_clk),
    .D(_00321_),
    .Q(\top_inst.grid_inst.data_path_wires[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _23789_ (.CLK(clknet_leaf_70_clk),
    .D(_00322_),
    .Q(\top_inst.grid_inst.data_path_wires[1][3] ));
 sky130_fd_sc_hd__dfxtp_4 _23790_ (.CLK(clknet_leaf_70_clk),
    .D(_00323_),
    .Q(\top_inst.grid_inst.data_path_wires[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _23791_ (.CLK(clknet_leaf_71_clk),
    .D(_00324_),
    .Q(\top_inst.grid_inst.data_path_wires[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _23792_ (.CLK(clknet_leaf_71_clk),
    .D(_00325_),
    .Q(\top_inst.grid_inst.data_path_wires[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _23793_ (.CLK(clknet_leaf_71_clk),
    .D(_00326_),
    .Q(\top_inst.grid_inst.data_path_wires[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _23794_ (.CLK(clknet_leaf_69_clk),
    .D(_00327_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _23795_ (.CLK(clknet_leaf_69_clk),
    .D(_00328_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _23796_ (.CLK(clknet_leaf_69_clk),
    .D(_00329_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _23797_ (.CLK(clknet_leaf_70_clk),
    .D(_00330_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _23798_ (.CLK(clknet_leaf_70_clk),
    .D(_00331_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _23799_ (.CLK(clknet_leaf_70_clk),
    .D(_00332_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23800_ (.CLK(clknet_leaf_70_clk),
    .D(_00333_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _23801_ (.CLK(clknet_leaf_72_clk),
    .D(_00334_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _23802_ (.CLK(clknet_leaf_77_clk),
    .D(_00335_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[0] ));
 sky130_fd_sc_hd__dfxtp_1 _23803_ (.CLK(clknet_leaf_77_clk),
    .D(_00336_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[1] ));
 sky130_fd_sc_hd__dfxtp_1 _23804_ (.CLK(clknet_leaf_77_clk),
    .D(_00337_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _23805_ (.CLK(clknet_leaf_69_clk),
    .D(_00338_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[3] ));
 sky130_fd_sc_hd__dfxtp_2 _23806_ (.CLK(clknet_leaf_76_clk),
    .D(_00339_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[4] ));
 sky130_fd_sc_hd__dfxtp_1 _23807_ (.CLK(clknet_leaf_74_clk),
    .D(_00340_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23808_ (.CLK(clknet_leaf_74_clk),
    .D(_00341_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[6] ));
 sky130_fd_sc_hd__dfxtp_1 _23809_ (.CLK(clknet_leaf_74_clk),
    .D(_00342_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[7] ));
 sky130_fd_sc_hd__dfxtp_1 _23810_ (.CLK(clknet_leaf_72_clk),
    .D(_00343_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[8] ));
 sky130_fd_sc_hd__dfxtp_1 _23811_ (.CLK(clknet_leaf_72_clk),
    .D(_00344_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[9] ));
 sky130_fd_sc_hd__dfxtp_1 _23812_ (.CLK(clknet_leaf_72_clk),
    .D(_00345_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[10] ));
 sky130_fd_sc_hd__dfxtp_1 _23813_ (.CLK(clknet_leaf_72_clk),
    .D(_00346_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[11] ));
 sky130_fd_sc_hd__dfxtp_1 _23814_ (.CLK(clknet_leaf_72_clk),
    .D(_00347_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[12] ));
 sky130_fd_sc_hd__dfxtp_1 _23815_ (.CLK(clknet_leaf_72_clk),
    .D(_00348_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _23816_ (.CLK(clknet_leaf_73_clk),
    .D(_00349_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[14] ));
 sky130_fd_sc_hd__dfxtp_1 _23817_ (.CLK(clknet_leaf_73_clk),
    .D(_00350_),
    .Q(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[15] ));
 sky130_fd_sc_hd__dfxtp_1 _23818_ (.CLK(clknet_leaf_93_clk),
    .D(_00351_),
    .Q(\top_inst.grid_inst.data_path_wires[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _23819_ (.CLK(clknet_leaf_93_clk),
    .D(_00352_),
    .Q(\top_inst.grid_inst.data_path_wires[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _23820_ (.CLK(clknet_leaf_93_clk),
    .D(_00353_),
    .Q(\top_inst.grid_inst.data_path_wires[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _23821_ (.CLK(clknet_leaf_93_clk),
    .D(_00354_),
    .Q(\top_inst.grid_inst.data_path_wires[2][3] ));
 sky130_fd_sc_hd__dfxtp_4 _23822_ (.CLK(clknet_leaf_93_clk),
    .D(_00355_),
    .Q(\top_inst.grid_inst.data_path_wires[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _23823_ (.CLK(clknet_leaf_94_clk),
    .D(_00356_),
    .Q(\top_inst.grid_inst.data_path_wires[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _23824_ (.CLK(clknet_leaf_94_clk),
    .D(_00357_),
    .Q(\top_inst.grid_inst.data_path_wires[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _23825_ (.CLK(clknet_leaf_94_clk),
    .D(_00358_),
    .Q(\top_inst.grid_inst.data_path_wires[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _23826_ (.CLK(clknet_leaf_93_clk),
    .D(_00359_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _23827_ (.CLK(clknet_leaf_93_clk),
    .D(_00360_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _23828_ (.CLK(clknet_leaf_93_clk),
    .D(_00361_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _23829_ (.CLK(clknet_leaf_93_clk),
    .D(_00362_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _23830_ (.CLK(clknet_leaf_94_clk),
    .D(_00363_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _23831_ (.CLK(clknet_leaf_93_clk),
    .D(_00364_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23832_ (.CLK(clknet_leaf_93_clk),
    .D(_00365_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _23833_ (.CLK(clknet_leaf_93_clk),
    .D(_00366_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _23834_ (.CLK(clknet_leaf_92_clk),
    .D(_00367_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[0] ));
 sky130_fd_sc_hd__dfxtp_1 _23835_ (.CLK(clknet_leaf_92_clk),
    .D(_00368_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[1] ));
 sky130_fd_sc_hd__dfxtp_1 _23836_ (.CLK(clknet_leaf_92_clk),
    .D(_00369_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _23837_ (.CLK(clknet_leaf_92_clk),
    .D(_00370_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[3] ));
 sky130_fd_sc_hd__dfxtp_1 _23838_ (.CLK(clknet_leaf_89_clk),
    .D(_00371_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[4] ));
 sky130_fd_sc_hd__dfxtp_1 _23839_ (.CLK(clknet_leaf_89_clk),
    .D(_00372_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23840_ (.CLK(clknet_leaf_89_clk),
    .D(_00373_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[6] ));
 sky130_fd_sc_hd__dfxtp_1 _23841_ (.CLK(clknet_leaf_96_clk),
    .D(_00374_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[7] ));
 sky130_fd_sc_hd__dfxtp_1 _23842_ (.CLK(clknet_leaf_96_clk),
    .D(_00375_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[8] ));
 sky130_fd_sc_hd__dfxtp_1 _23843_ (.CLK(clknet_leaf_96_clk),
    .D(_00376_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[9] ));
 sky130_fd_sc_hd__dfxtp_1 _23844_ (.CLK(clknet_leaf_96_clk),
    .D(_00377_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[10] ));
 sky130_fd_sc_hd__dfxtp_1 _23845_ (.CLK(clknet_leaf_96_clk),
    .D(_00378_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[11] ));
 sky130_fd_sc_hd__dfxtp_1 _23846_ (.CLK(clknet_leaf_95_clk),
    .D(_00379_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[12] ));
 sky130_fd_sc_hd__dfxtp_1 _23847_ (.CLK(clknet_leaf_95_clk),
    .D(_00380_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _23848_ (.CLK(clknet_leaf_95_clk),
    .D(_00381_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[14] ));
 sky130_fd_sc_hd__dfxtp_1 _23849_ (.CLK(clknet_leaf_95_clk),
    .D(_00382_),
    .Q(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[15] ));
 sky130_fd_sc_hd__dfxtp_2 _23850_ (.CLK(clknet_leaf_68_clk),
    .D(_00383_),
    .Q(\top_inst.grid_inst.data_path_wires[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _23851_ (.CLK(clknet_leaf_68_clk),
    .D(_00384_),
    .Q(\top_inst.grid_inst.data_path_wires[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _23852_ (.CLK(clknet_leaf_68_clk),
    .D(_00385_),
    .Q(\top_inst.grid_inst.data_path_wires[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _23853_ (.CLK(clknet_leaf_68_clk),
    .D(_00386_),
    .Q(\top_inst.grid_inst.data_path_wires[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _23854_ (.CLK(clknet_leaf_69_clk),
    .D(_00387_),
    .Q(\top_inst.grid_inst.data_path_wires[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _23855_ (.CLK(clknet_leaf_70_clk),
    .D(_00388_),
    .Q(\top_inst.grid_inst.data_path_wires[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _23856_ (.CLK(clknet_leaf_69_clk),
    .D(_00389_),
    .Q(\top_inst.grid_inst.data_path_wires[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 _23857_ (.CLK(clknet_leaf_68_clk),
    .D(_00390_),
    .Q(\top_inst.grid_inst.data_path_wires[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _23858_ (.CLK(clknet_leaf_77_clk),
    .D(_00391_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _23859_ (.CLK(clknet_leaf_77_clk),
    .D(_00392_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _23860_ (.CLK(clknet_leaf_77_clk),
    .D(_00393_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _23861_ (.CLK(clknet_leaf_77_clk),
    .D(_00394_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _23862_ (.CLK(clknet_leaf_68_clk),
    .D(_00395_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _23863_ (.CLK(clknet_leaf_68_clk),
    .D(_00396_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23864_ (.CLK(clknet_leaf_68_clk),
    .D(_00397_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _23865_ (.CLK(clknet_leaf_68_clk),
    .D(_00398_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _23866_ (.CLK(clknet_leaf_78_clk),
    .D(_00399_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[0] ));
 sky130_fd_sc_hd__dfxtp_1 _23867_ (.CLK(clknet_leaf_78_clk),
    .D(_00400_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[1] ));
 sky130_fd_sc_hd__dfxtp_2 _23868_ (.CLK(clknet_leaf_78_clk),
    .D(_00401_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _23869_ (.CLK(clknet_leaf_78_clk),
    .D(_00402_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[3] ));
 sky130_fd_sc_hd__dfxtp_1 _23870_ (.CLK(clknet_leaf_78_clk),
    .D(_00403_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[4] ));
 sky130_fd_sc_hd__dfxtp_1 _23871_ (.CLK(clknet_leaf_78_clk),
    .D(_00404_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23872_ (.CLK(clknet_leaf_78_clk),
    .D(_00405_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[6] ));
 sky130_fd_sc_hd__dfxtp_1 _23873_ (.CLK(clknet_leaf_50_clk),
    .D(_00406_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[7] ));
 sky130_fd_sc_hd__dfxtp_1 _23874_ (.CLK(clknet_leaf_50_clk),
    .D(_00407_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[8] ));
 sky130_fd_sc_hd__dfxtp_1 _23875_ (.CLK(clknet_leaf_51_clk),
    .D(_00408_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[9] ));
 sky130_fd_sc_hd__dfxtp_1 _23876_ (.CLK(clknet_leaf_62_clk),
    .D(_00409_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[10] ));
 sky130_fd_sc_hd__dfxtp_1 _23877_ (.CLK(clknet_leaf_51_clk),
    .D(_00410_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[11] ));
 sky130_fd_sc_hd__dfxtp_1 _23878_ (.CLK(clknet_leaf_51_clk),
    .D(_00411_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[12] ));
 sky130_fd_sc_hd__dfxtp_1 _23879_ (.CLK(clknet_leaf_61_clk),
    .D(_00412_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _23880_ (.CLK(clknet_leaf_62_clk),
    .D(_00413_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[14] ));
 sky130_fd_sc_hd__dfxtp_1 _23881_ (.CLK(clknet_leaf_50_clk),
    .D(_00414_),
    .Q(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[15] ));
 sky130_fd_sc_hd__dfxtp_2 _23882_ (.CLK(clknet_leaf_63_clk),
    .D(_00415_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _23883_ (.CLK(clknet_leaf_61_clk),
    .D(_00416_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _23884_ (.CLK(clknet_leaf_61_clk),
    .D(_00417_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_4 _23885_ (.CLK(clknet_leaf_64_clk),
    .D(_00418_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_4 _23886_ (.CLK(clknet_leaf_64_clk),
    .D(_00419_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _23887_ (.CLK(clknet_leaf_64_clk),
    .D(_00420_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23888_ (.CLK(clknet_leaf_64_clk),
    .D(_00421_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _23889_ (.CLK(clknet_leaf_63_clk),
    .D(_00422_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _23890_ (.CLK(clknet_leaf_62_clk),
    .D(_00423_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[0] ));
 sky130_fd_sc_hd__dfxtp_1 _23891_ (.CLK(clknet_leaf_51_clk),
    .D(_00424_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[1] ));
 sky130_fd_sc_hd__dfxtp_1 _23892_ (.CLK(clknet_leaf_62_clk),
    .D(_00425_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _23893_ (.CLK(clknet_leaf_52_clk),
    .D(_00426_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[3] ));
 sky130_fd_sc_hd__dfxtp_1 _23894_ (.CLK(clknet_leaf_51_clk),
    .D(_00427_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[4] ));
 sky130_fd_sc_hd__dfxtp_1 _23895_ (.CLK(clknet_leaf_51_clk),
    .D(_00428_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23896_ (.CLK(clknet_leaf_52_clk),
    .D(_00429_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[6] ));
 sky130_fd_sc_hd__dfxtp_1 _23897_ (.CLK(clknet_leaf_52_clk),
    .D(_00430_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[7] ));
 sky130_fd_sc_hd__dfxtp_1 _23898_ (.CLK(clknet_leaf_52_clk),
    .D(_00431_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[8] ));
 sky130_fd_sc_hd__dfxtp_1 _23899_ (.CLK(clknet_leaf_52_clk),
    .D(_00432_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[9] ));
 sky130_fd_sc_hd__dfxtp_2 _23900_ (.CLK(clknet_leaf_51_clk),
    .D(_00433_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[10] ));
 sky130_fd_sc_hd__dfxtp_2 _23901_ (.CLK(clknet_4_13__leaf_clk),
    .D(_00434_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[11] ));
 sky130_fd_sc_hd__dfxtp_2 _23902_ (.CLK(clknet_leaf_52_clk),
    .D(_00435_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[12] ));
 sky130_fd_sc_hd__dfxtp_2 _23903_ (.CLK(clknet_leaf_59_clk),
    .D(_00436_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[13] ));
 sky130_fd_sc_hd__dfxtp_2 _23904_ (.CLK(clknet_leaf_52_clk),
    .D(_00437_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[14] ));
 sky130_fd_sc_hd__dfxtp_2 _23905_ (.CLK(clknet_leaf_54_clk),
    .D(_00438_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[15] ));
 sky130_fd_sc_hd__dfxtp_1 _23906_ (.CLK(clknet_leaf_37_clk),
    .D(_00439_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[16] ));
 sky130_fd_sc_hd__dfxtp_1 _23907_ (.CLK(clknet_leaf_37_clk),
    .D(_00440_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[17] ));
 sky130_fd_sc_hd__dfxtp_1 _23908_ (.CLK(clknet_leaf_36_clk),
    .D(_00441_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[18] ));
 sky130_fd_sc_hd__dfxtp_1 _23909_ (.CLK(clknet_leaf_36_clk),
    .D(_00442_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[19] ));
 sky130_fd_sc_hd__dfxtp_1 _23910_ (.CLK(clknet_leaf_36_clk),
    .D(_00443_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[20] ));
 sky130_fd_sc_hd__dfxtp_1 _23911_ (.CLK(clknet_leaf_36_clk),
    .D(_00444_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[21] ));
 sky130_fd_sc_hd__dfxtp_1 _23912_ (.CLK(clknet_leaf_33_clk),
    .D(_00445_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[23] ));
 sky130_fd_sc_hd__dfxtp_1 _23913_ (.CLK(clknet_leaf_33_clk),
    .D(_00446_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[24] ));
 sky130_fd_sc_hd__dfxtp_2 _23914_ (.CLK(clknet_leaf_35_clk),
    .D(_00447_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[25] ));
 sky130_fd_sc_hd__dfxtp_1 _23915_ (.CLK(clknet_leaf_33_clk),
    .D(_00448_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[27] ));
 sky130_fd_sc_hd__dfxtp_1 _23916_ (.CLK(clknet_leaf_35_clk),
    .D(_00449_),
    .Q(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[31] ));
 sky130_fd_sc_hd__dfxtp_2 _23917_ (.CLK(clknet_leaf_77_clk),
    .D(_00450_),
    .Q(\top_inst.grid_inst.data_path_wires[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _23918_ (.CLK(clknet_leaf_77_clk),
    .D(_00451_),
    .Q(\top_inst.grid_inst.data_path_wires[6][1] ));
 sky130_fd_sc_hd__dfxtp_2 _23919_ (.CLK(clknet_leaf_77_clk),
    .D(_00452_),
    .Q(\top_inst.grid_inst.data_path_wires[6][2] ));
 sky130_fd_sc_hd__dfxtp_4 _23920_ (.CLK(clknet_leaf_76_clk),
    .D(_00453_),
    .Q(\top_inst.grid_inst.data_path_wires[6][3] ));
 sky130_fd_sc_hd__dfxtp_2 _23921_ (.CLK(clknet_leaf_77_clk),
    .D(_00454_),
    .Q(\top_inst.grid_inst.data_path_wires[6][4] ));
 sky130_fd_sc_hd__dfxtp_2 _23922_ (.CLK(clknet_leaf_77_clk),
    .D(_00455_),
    .Q(\top_inst.grid_inst.data_path_wires[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _23923_ (.CLK(clknet_leaf_76_clk),
    .D(_00456_),
    .Q(\top_inst.grid_inst.data_path_wires[6][6] ));
 sky130_fd_sc_hd__dfxtp_2 _23924_ (.CLK(clknet_leaf_76_clk),
    .D(_00457_),
    .Q(\top_inst.grid_inst.data_path_wires[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _23925_ (.CLK(clknet_leaf_76_clk),
    .D(_00458_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _23926_ (.CLK(clknet_leaf_76_clk),
    .D(_00459_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _23927_ (.CLK(clknet_leaf_76_clk),
    .D(_00460_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_4 _23928_ (.CLK(clknet_leaf_76_clk),
    .D(_00461_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_4 _23929_ (.CLK(clknet_leaf_76_clk),
    .D(_00462_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _23930_ (.CLK(clknet_leaf_75_clk),
    .D(_00463_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23931_ (.CLK(clknet_leaf_75_clk),
    .D(_00464_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _23932_ (.CLK(clknet_leaf_91_clk),
    .D(_00465_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_2 _23933_ (.CLK(clknet_leaf_85_clk),
    .D(_00466_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[0] ));
 sky130_fd_sc_hd__dfxtp_1 _23934_ (.CLK(clknet_leaf_81_clk),
    .D(_00467_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[1] ));
 sky130_fd_sc_hd__dfxtp_2 _23935_ (.CLK(clknet_leaf_81_clk),
    .D(_00468_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _23936_ (.CLK(clknet_leaf_80_clk),
    .D(_00469_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[3] ));
 sky130_fd_sc_hd__dfxtp_2 _23937_ (.CLK(clknet_leaf_80_clk),
    .D(_00470_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[4] ));
 sky130_fd_sc_hd__dfxtp_2 _23938_ (.CLK(clknet_leaf_81_clk),
    .D(_00471_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23939_ (.CLK(clknet_leaf_81_clk),
    .D(_00472_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[6] ));
 sky130_fd_sc_hd__dfxtp_2 _23940_ (.CLK(clknet_leaf_81_clk),
    .D(_00473_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[7] ));
 sky130_fd_sc_hd__dfxtp_1 _23941_ (.CLK(clknet_leaf_81_clk),
    .D(_00474_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[8] ));
 sky130_fd_sc_hd__dfxtp_1 _23942_ (.CLK(clknet_leaf_81_clk),
    .D(_00475_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[9] ));
 sky130_fd_sc_hd__dfxtp_1 _23943_ (.CLK(clknet_leaf_85_clk),
    .D(_00476_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[10] ));
 sky130_fd_sc_hd__dfxtp_1 _23944_ (.CLK(clknet_leaf_91_clk),
    .D(_00477_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[11] ));
 sky130_fd_sc_hd__dfxtp_1 _23945_ (.CLK(clknet_leaf_85_clk),
    .D(_00478_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[12] ));
 sky130_fd_sc_hd__dfxtp_1 _23946_ (.CLK(clknet_leaf_90_clk),
    .D(_00479_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _23947_ (.CLK(clknet_leaf_85_clk),
    .D(_00480_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[14] ));
 sky130_fd_sc_hd__dfxtp_1 _23948_ (.CLK(clknet_leaf_81_clk),
    .D(_00481_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[15] ));
 sky130_fd_sc_hd__dfxtp_1 _23949_ (.CLK(clknet_leaf_81_clk),
    .D(_00482_),
    .Q(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[16] ));
 sky130_fd_sc_hd__dfxtp_2 _23950_ (.CLK(clknet_leaf_90_clk),
    .D(_00483_),
    .Q(\top_inst.grid_inst.data_path_wires[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _23951_ (.CLK(clknet_leaf_90_clk),
    .D(_00484_),
    .Q(\top_inst.grid_inst.data_path_wires[7][1] ));
 sky130_fd_sc_hd__dfxtp_2 _23952_ (.CLK(clknet_leaf_90_clk),
    .D(_00485_),
    .Q(\top_inst.grid_inst.data_path_wires[7][2] ));
 sky130_fd_sc_hd__dfxtp_2 _23953_ (.CLK(clknet_leaf_90_clk),
    .D(_00486_),
    .Q(\top_inst.grid_inst.data_path_wires[7][3] ));
 sky130_fd_sc_hd__dfxtp_2 _23954_ (.CLK(clknet_leaf_91_clk),
    .D(_00487_),
    .Q(\top_inst.grid_inst.data_path_wires[7][4] ));
 sky130_fd_sc_hd__dfxtp_2 _23955_ (.CLK(clknet_leaf_91_clk),
    .D(_00488_),
    .Q(\top_inst.grid_inst.data_path_wires[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _23956_ (.CLK(clknet_leaf_91_clk),
    .D(_00489_),
    .Q(\top_inst.grid_inst.data_path_wires[7][6] ));
 sky130_fd_sc_hd__dfxtp_4 _23957_ (.CLK(clknet_leaf_91_clk),
    .D(_00490_),
    .Q(\top_inst.grid_inst.data_path_wires[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _23958_ (.CLK(clknet_leaf_89_clk),
    .D(_00491_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _23959_ (.CLK(clknet_leaf_89_clk),
    .D(_00492_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _23960_ (.CLK(clknet_leaf_89_clk),
    .D(_00493_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _23961_ (.CLK(clknet_leaf_89_clk),
    .D(_00494_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _23962_ (.CLK(clknet_leaf_89_clk),
    .D(_00495_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _23963_ (.CLK(clknet_leaf_88_clk),
    .D(_00496_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23964_ (.CLK(clknet_leaf_88_clk),
    .D(_00497_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _23965_ (.CLK(clknet_leaf_89_clk),
    .D(_00498_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_2 _23966_ (.CLK(clknet_leaf_85_clk),
    .D(_00499_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[0] ));
 sky130_fd_sc_hd__dfxtp_2 _23967_ (.CLK(clknet_leaf_90_clk),
    .D(_00500_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[1] ));
 sky130_fd_sc_hd__dfxtp_2 _23968_ (.CLK(clknet_leaf_86_clk),
    .D(_00501_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[2] ));
 sky130_fd_sc_hd__dfxtp_2 _23969_ (.CLK(clknet_leaf_85_clk),
    .D(_00502_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[3] ));
 sky130_fd_sc_hd__dfxtp_2 _23970_ (.CLK(clknet_leaf_85_clk),
    .D(_00503_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[4] ));
 sky130_fd_sc_hd__dfxtp_2 _23971_ (.CLK(clknet_leaf_86_clk),
    .D(_00504_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23972_ (.CLK(clknet_leaf_114_clk),
    .D(_00505_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[6] ));
 sky130_fd_sc_hd__dfxtp_2 _23973_ (.CLK(clknet_leaf_86_clk),
    .D(_00506_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[7] ));
 sky130_fd_sc_hd__dfxtp_2 _23974_ (.CLK(clknet_leaf_87_clk),
    .D(_00507_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[8] ));
 sky130_fd_sc_hd__dfxtp_2 _23975_ (.CLK(clknet_leaf_87_clk),
    .D(_00508_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[9] ));
 sky130_fd_sc_hd__dfxtp_2 _23976_ (.CLK(clknet_leaf_87_clk),
    .D(_00509_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[10] ));
 sky130_fd_sc_hd__dfxtp_2 _23977_ (.CLK(clknet_leaf_87_clk),
    .D(_00510_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[11] ));
 sky130_fd_sc_hd__dfxtp_2 _23978_ (.CLK(clknet_leaf_87_clk),
    .D(_00511_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[12] ));
 sky130_fd_sc_hd__dfxtp_1 _23979_ (.CLK(clknet_leaf_87_clk),
    .D(_00512_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _23980_ (.CLK(clknet_leaf_87_clk),
    .D(_00513_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[14] ));
 sky130_fd_sc_hd__dfxtp_2 _23981_ (.CLK(clknet_leaf_88_clk),
    .D(_00514_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[15] ));
 sky130_fd_sc_hd__dfxtp_2 _23982_ (.CLK(clknet_leaf_87_clk),
    .D(_00515_),
    .Q(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[16] ));
 sky130_fd_sc_hd__dfxtp_2 _23983_ (.CLK(clknet_leaf_81_clk),
    .D(_00516_),
    .Q(\top_inst.grid_inst.data_path_wires[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 _23984_ (.CLK(clknet_leaf_80_clk),
    .D(_00517_),
    .Q(\top_inst.grid_inst.data_path_wires[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _23985_ (.CLK(clknet_leaf_80_clk),
    .D(_00518_),
    .Q(\top_inst.grid_inst.data_path_wires[8][2] ));
 sky130_fd_sc_hd__dfxtp_2 _23986_ (.CLK(clknet_leaf_80_clk),
    .D(_00519_),
    .Q(\top_inst.grid_inst.data_path_wires[8][3] ));
 sky130_fd_sc_hd__dfxtp_2 _23987_ (.CLK(clknet_leaf_80_clk),
    .D(_00520_),
    .Q(\top_inst.grid_inst.data_path_wires[8][4] ));
 sky130_fd_sc_hd__dfxtp_2 _23988_ (.CLK(clknet_leaf_80_clk),
    .D(_00521_),
    .Q(\top_inst.grid_inst.data_path_wires[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _23989_ (.CLK(clknet_leaf_78_clk),
    .D(_00522_),
    .Q(\top_inst.grid_inst.data_path_wires[8][6] ));
 sky130_fd_sc_hd__dfxtp_2 _23990_ (.CLK(clknet_leaf_78_clk),
    .D(_00523_),
    .Q(\top_inst.grid_inst.data_path_wires[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _23991_ (.CLK(clknet_leaf_79_clk),
    .D(_00524_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _23992_ (.CLK(clknet_leaf_79_clk),
    .D(_00525_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _23993_ (.CLK(clknet_leaf_79_clk),
    .D(_00526_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _23994_ (.CLK(clknet_leaf_82_clk),
    .D(_00527_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _23995_ (.CLK(clknet_leaf_79_clk),
    .D(_00528_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _23996_ (.CLK(clknet_4_14__leaf_clk),
    .D(_00529_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _23997_ (.CLK(clknet_leaf_79_clk),
    .D(_00530_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _23998_ (.CLK(clknet_leaf_79_clk),
    .D(_00531_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_2 _23999_ (.CLK(clknet_leaf_81_clk),
    .D(net1069),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[0] ));
 sky130_fd_sc_hd__dfxtp_2 _24000_ (.CLK(clknet_leaf_83_clk),
    .D(_00533_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[1] ));
 sky130_fd_sc_hd__dfxtp_2 _24001_ (.CLK(clknet_leaf_81_clk),
    .D(_00534_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[2] ));
 sky130_fd_sc_hd__dfxtp_2 _24002_ (.CLK(clknet_leaf_46_clk),
    .D(_00535_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[3] ));
 sky130_fd_sc_hd__dfxtp_4 _24003_ (.CLK(clknet_leaf_82_clk),
    .D(_00536_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[4] ));
 sky130_fd_sc_hd__dfxtp_2 _24004_ (.CLK(clknet_leaf_82_clk),
    .D(_00537_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[5] ));
 sky130_fd_sc_hd__dfxtp_2 _24005_ (.CLK(clknet_leaf_46_clk),
    .D(_00538_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[6] ));
 sky130_fd_sc_hd__dfxtp_2 _24006_ (.CLK(clknet_leaf_46_clk),
    .D(_00539_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[7] ));
 sky130_fd_sc_hd__dfxtp_2 _24007_ (.CLK(clknet_leaf_46_clk),
    .D(_00540_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[8] ));
 sky130_fd_sc_hd__dfxtp_2 _24008_ (.CLK(clknet_leaf_47_clk),
    .D(_00541_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[9] ));
 sky130_fd_sc_hd__dfxtp_2 _24009_ (.CLK(clknet_leaf_47_clk),
    .D(_00542_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[10] ));
 sky130_fd_sc_hd__dfxtp_2 _24010_ (.CLK(clknet_leaf_47_clk),
    .D(_00543_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[11] ));
 sky130_fd_sc_hd__dfxtp_2 _24011_ (.CLK(clknet_leaf_47_clk),
    .D(_00544_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[12] ));
 sky130_fd_sc_hd__dfxtp_2 _24012_ (.CLK(clknet_leaf_47_clk),
    .D(_00545_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[13] ));
 sky130_fd_sc_hd__dfxtp_2 _24013_ (.CLK(clknet_leaf_48_clk),
    .D(_00546_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[14] ));
 sky130_fd_sc_hd__dfxtp_2 _24014_ (.CLK(clknet_leaf_48_clk),
    .D(_00547_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[15] ));
 sky130_fd_sc_hd__dfxtp_2 _24015_ (.CLK(clknet_leaf_48_clk),
    .D(_00548_),
    .Q(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[16] ));
 sky130_fd_sc_hd__dfxtp_1 _24016_ (.CLK(clknet_leaf_52_clk),
    .D(_00549_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _24017_ (.CLK(clknet_leaf_52_clk),
    .D(_00550_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _24018_ (.CLK(clknet_leaf_54_clk),
    .D(_00551_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _24019_ (.CLK(clknet_leaf_54_clk),
    .D(_00552_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_4 _24020_ (.CLK(clknet_leaf_54_clk),
    .D(_00553_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24021_ (.CLK(clknet_leaf_55_clk),
    .D(_00554_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _24022_ (.CLK(clknet_leaf_55_clk),
    .D(_00555_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24023_ (.CLK(clknet_leaf_53_clk),
    .D(_00556_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24024_ (.CLK(clknet_leaf_48_clk),
    .D(_00557_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[0] ));
 sky130_fd_sc_hd__dfxtp_1 _24025_ (.CLK(clknet_4_12__leaf_clk),
    .D(_00558_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24026_ (.CLK(clknet_leaf_48_clk),
    .D(_00559_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _24027_ (.CLK(clknet_leaf_48_clk),
    .D(_00560_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[3] ));
 sky130_fd_sc_hd__dfxtp_1 _24028_ (.CLK(clknet_leaf_48_clk),
    .D(_00561_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24029_ (.CLK(clknet_leaf_48_clk),
    .D(_00562_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[5] ));
 sky130_fd_sc_hd__dfxtp_1 _24030_ (.CLK(clknet_leaf_41_clk),
    .D(_00563_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24031_ (.CLK(clknet_leaf_48_clk),
    .D(_00564_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24032_ (.CLK(clknet_leaf_53_clk),
    .D(_00565_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[8] ));
 sky130_fd_sc_hd__dfxtp_1 _24033_ (.CLK(clknet_leaf_41_clk),
    .D(_00566_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[9] ));
 sky130_fd_sc_hd__dfxtp_1 _24034_ (.CLK(clknet_leaf_41_clk),
    .D(_00567_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[10] ));
 sky130_fd_sc_hd__dfxtp_1 _24035_ (.CLK(clknet_leaf_41_clk),
    .D(_00568_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[11] ));
 sky130_fd_sc_hd__dfxtp_1 _24036_ (.CLK(clknet_leaf_41_clk),
    .D(_00569_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[12] ));
 sky130_fd_sc_hd__dfxtp_1 _24037_ (.CLK(clknet_leaf_42_clk),
    .D(_00570_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _24038_ (.CLK(clknet_leaf_42_clk),
    .D(_00571_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[14] ));
 sky130_fd_sc_hd__dfxtp_1 _24039_ (.CLK(clknet_leaf_42_clk),
    .D(_00572_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[15] ));
 sky130_fd_sc_hd__dfxtp_1 _24040_ (.CLK(clknet_leaf_42_clk),
    .D(_00573_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[16] ));
 sky130_fd_sc_hd__dfxtp_1 _24041_ (.CLK(clknet_leaf_42_clk),
    .D(_00574_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[17] ));
 sky130_fd_sc_hd__dfxtp_1 _24042_ (.CLK(clknet_leaf_42_clk),
    .D(_00575_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[18] ));
 sky130_fd_sc_hd__dfxtp_1 _24043_ (.CLK(clknet_leaf_42_clk),
    .D(_00576_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[19] ));
 sky130_fd_sc_hd__dfxtp_1 _24044_ (.CLK(clknet_leaf_42_clk),
    .D(_00577_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[20] ));
 sky130_fd_sc_hd__dfxtp_1 _24045_ (.CLK(clknet_leaf_42_clk),
    .D(_00578_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[21] ));
 sky130_fd_sc_hd__dfxtp_1 _24046_ (.CLK(clknet_4_7__leaf_clk),
    .D(_00579_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[22] ));
 sky130_fd_sc_hd__dfxtp_1 _24047_ (.CLK(clknet_leaf_34_clk),
    .D(_00580_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[23] ));
 sky130_fd_sc_hd__dfxtp_1 _24048_ (.CLK(clknet_leaf_34_clk),
    .D(_00581_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[24] ));
 sky130_fd_sc_hd__dfxtp_1 _24049_ (.CLK(clknet_leaf_34_clk),
    .D(_00582_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[25] ));
 sky130_fd_sc_hd__dfxtp_1 _24050_ (.CLK(clknet_leaf_34_clk),
    .D(_00583_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[26] ));
 sky130_fd_sc_hd__dfxtp_1 _24051_ (.CLK(clknet_leaf_34_clk),
    .D(_00584_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[27] ));
 sky130_fd_sc_hd__dfxtp_1 _24052_ (.CLK(clknet_leaf_34_clk),
    .D(_00585_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[28] ));
 sky130_fd_sc_hd__dfxtp_1 _24053_ (.CLK(clknet_leaf_34_clk),
    .D(_00586_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[29] ));
 sky130_fd_sc_hd__dfxtp_1 _24054_ (.CLK(clknet_leaf_34_clk),
    .D(_00587_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[30] ));
 sky130_fd_sc_hd__dfxtp_1 _24055_ (.CLK(clknet_leaf_34_clk),
    .D(_00588_),
    .Q(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[31] ));
 sky130_fd_sc_hd__dfxtp_2 _24056_ (.CLK(clknet_leaf_46_clk),
    .D(_00589_),
    .Q(\top_inst.grid_inst.data_path_wires[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _24057_ (.CLK(clknet_leaf_46_clk),
    .D(_00590_),
    .Q(\top_inst.grid_inst.data_path_wires[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 _24058_ (.CLK(clknet_leaf_83_clk),
    .D(_00591_),
    .Q(\top_inst.grid_inst.data_path_wires[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 _24059_ (.CLK(clknet_leaf_45_clk),
    .D(_00592_),
    .Q(\top_inst.grid_inst.data_path_wires[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 _24060_ (.CLK(clknet_leaf_45_clk),
    .D(_00593_),
    .Q(\top_inst.grid_inst.data_path_wires[11][4] ));
 sky130_fd_sc_hd__dfxtp_2 _24061_ (.CLK(clknet_leaf_45_clk),
    .D(_00594_),
    .Q(\top_inst.grid_inst.data_path_wires[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _24062_ (.CLK(clknet_leaf_84_clk),
    .D(_00595_),
    .Q(\top_inst.grid_inst.data_path_wires[11][6] ));
 sky130_fd_sc_hd__dfxtp_2 _24063_ (.CLK(clknet_leaf_83_clk),
    .D(_00596_),
    .Q(\top_inst.grid_inst.data_path_wires[11][7] ));
 sky130_fd_sc_hd__dfxtp_2 _24064_ (.CLK(clknet_leaf_83_clk),
    .D(_00597_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _24065_ (.CLK(clknet_leaf_83_clk),
    .D(_00598_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24066_ (.CLK(clknet_leaf_84_clk),
    .D(_00599_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _24067_ (.CLK(clknet_leaf_84_clk),
    .D(_00600_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _24068_ (.CLK(clknet_leaf_84_clk),
    .D(_00601_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24069_ (.CLK(clknet_leaf_84_clk),
    .D(_00602_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _24070_ (.CLK(clknet_leaf_84_clk),
    .D(_00603_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24071_ (.CLK(clknet_leaf_84_clk),
    .D(_00604_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24072_ (.CLK(clknet_leaf_114_clk),
    .D(_00605_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[0] ));
 sky130_fd_sc_hd__dfxtp_1 _24073_ (.CLK(clknet_leaf_114_clk),
    .D(_00606_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24074_ (.CLK(clknet_leaf_112_clk),
    .D(_00607_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _24075_ (.CLK(clknet_leaf_114_clk),
    .D(_00608_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[3] ));
 sky130_fd_sc_hd__dfxtp_1 _24076_ (.CLK(clknet_leaf_112_clk),
    .D(_00609_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24077_ (.CLK(clknet_leaf_113_clk),
    .D(_00610_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[5] ));
 sky130_fd_sc_hd__dfxtp_1 _24078_ (.CLK(clknet_leaf_113_clk),
    .D(_00611_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24079_ (.CLK(clknet_leaf_113_clk),
    .D(_00612_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24080_ (.CLK(clknet_leaf_113_clk),
    .D(_00613_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[8] ));
 sky130_fd_sc_hd__dfxtp_1 _24081_ (.CLK(clknet_leaf_111_clk),
    .D(_00614_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[9] ));
 sky130_fd_sc_hd__dfxtp_1 _24082_ (.CLK(clknet_leaf_111_clk),
    .D(_00615_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[10] ));
 sky130_fd_sc_hd__dfxtp_1 _24083_ (.CLK(clknet_leaf_87_clk),
    .D(_00616_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[11] ));
 sky130_fd_sc_hd__dfxtp_1 _24084_ (.CLK(clknet_leaf_87_clk),
    .D(_00617_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[12] ));
 sky130_fd_sc_hd__dfxtp_1 _24085_ (.CLK(clknet_leaf_87_clk),
    .D(_00618_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _24086_ (.CLK(clknet_leaf_87_clk),
    .D(_00619_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[14] ));
 sky130_fd_sc_hd__dfxtp_1 _24087_ (.CLK(clknet_leaf_86_clk),
    .D(_00620_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[15] ));
 sky130_fd_sc_hd__dfxtp_1 _24088_ (.CLK(clknet_leaf_87_clk),
    .D(_00621_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[16] ));
 sky130_fd_sc_hd__dfxtp_1 _24089_ (.CLK(clknet_leaf_97_clk),
    .D(_00622_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[17] ));
 sky130_fd_sc_hd__dfxtp_1 _24090_ (.CLK(clknet_leaf_97_clk),
    .D(_00623_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[18] ));
 sky130_fd_sc_hd__dfxtp_1 _24091_ (.CLK(clknet_leaf_97_clk),
    .D(_00624_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[19] ));
 sky130_fd_sc_hd__dfxtp_1 _24092_ (.CLK(clknet_leaf_99_clk),
    .D(_00625_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[20] ));
 sky130_fd_sc_hd__dfxtp_1 _24093_ (.CLK(clknet_leaf_99_clk),
    .D(_00626_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[21] ));
 sky130_fd_sc_hd__dfxtp_1 _24094_ (.CLK(clknet_leaf_99_clk),
    .D(_00627_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[23] ));
 sky130_fd_sc_hd__dfxtp_1 _24095_ (.CLK(clknet_leaf_99_clk),
    .D(_00628_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[24] ));
 sky130_fd_sc_hd__dfxtp_1 _24096_ (.CLK(clknet_leaf_99_clk),
    .D(_00629_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[25] ));
 sky130_fd_sc_hd__dfxtp_1 _24097_ (.CLK(clknet_leaf_99_clk),
    .D(_00630_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[27] ));
 sky130_fd_sc_hd__dfxtp_1 _24098_ (.CLK(clknet_leaf_97_clk),
    .D(_00631_),
    .Q(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[31] ));
 sky130_fd_sc_hd__dfxtp_1 _24099_ (.CLK(clknet_leaf_15_clk),
    .D(_00632_),
    .Q(\top_inst.grid_inst.data_path_wires[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 _24100_ (.CLK(clknet_leaf_15_clk),
    .D(_00633_),
    .Q(\top_inst.grid_inst.data_path_wires[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _24101_ (.CLK(clknet_leaf_15_clk),
    .D(_00634_),
    .Q(\top_inst.grid_inst.data_path_wires[12][2] ));
 sky130_fd_sc_hd__dfxtp_2 _24102_ (.CLK(clknet_leaf_15_clk),
    .D(_00635_),
    .Q(\top_inst.grid_inst.data_path_wires[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 _24103_ (.CLK(clknet_leaf_115_clk),
    .D(_00636_),
    .Q(\top_inst.grid_inst.data_path_wires[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 _24104_ (.CLK(clknet_leaf_15_clk),
    .D(_00637_),
    .Q(\top_inst.grid_inst.data_path_wires[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _24105_ (.CLK(clknet_leaf_15_clk),
    .D(_00638_),
    .Q(\top_inst.grid_inst.data_path_wires[12][6] ));
 sky130_fd_sc_hd__dfxtp_2 _24106_ (.CLK(clknet_leaf_115_clk),
    .D(_00639_),
    .Q(\top_inst.grid_inst.data_path_wires[12][7] ));
 sky130_fd_sc_hd__dfxtp_2 _24107_ (.CLK(clknet_leaf_14_clk),
    .D(_00640_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _24108_ (.CLK(clknet_leaf_14_clk),
    .D(_00641_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24109_ (.CLK(clknet_leaf_16_clk),
    .D(_00642_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _24110_ (.CLK(clknet_leaf_14_clk),
    .D(_00643_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _24111_ (.CLK(clknet_leaf_16_clk),
    .D(_00644_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24112_ (.CLK(clknet_leaf_16_clk),
    .D(_00645_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _24113_ (.CLK(clknet_leaf_16_clk),
    .D(_00646_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24114_ (.CLK(clknet_leaf_16_clk),
    .D(_00647_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24115_ (.CLK(clknet_leaf_118_clk),
    .D(_00648_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[0] ));
 sky130_fd_sc_hd__dfxtp_1 _24116_ (.CLK(clknet_leaf_12_clk),
    .D(_00649_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24117_ (.CLK(clknet_leaf_12_clk),
    .D(_00650_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _24118_ (.CLK(clknet_leaf_13_clk),
    .D(_00651_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[3] ));
 sky130_fd_sc_hd__dfxtp_1 _24119_ (.CLK(clknet_leaf_13_clk),
    .D(_00652_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24120_ (.CLK(clknet_leaf_13_clk),
    .D(_00653_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[5] ));
 sky130_fd_sc_hd__dfxtp_1 _24121_ (.CLK(clknet_leaf_13_clk),
    .D(_00654_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24122_ (.CLK(clknet_leaf_12_clk),
    .D(_00655_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[7] ));
 sky130_fd_sc_hd__dfxtp_2 _24123_ (.CLK(clknet_leaf_11_clk),
    .D(_00656_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[8] ));
 sky130_fd_sc_hd__dfxtp_1 _24124_ (.CLK(clknet_leaf_118_clk),
    .D(_00657_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[9] ));
 sky130_fd_sc_hd__dfxtp_2 _24125_ (.CLK(clknet_leaf_119_clk),
    .D(_00658_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[10] ));
 sky130_fd_sc_hd__dfxtp_1 _24126_ (.CLK(clknet_leaf_118_clk),
    .D(_00659_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[11] ));
 sky130_fd_sc_hd__dfxtp_1 _24127_ (.CLK(clknet_leaf_118_clk),
    .D(_00660_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[12] ));
 sky130_fd_sc_hd__dfxtp_2 _24128_ (.CLK(clknet_leaf_117_clk),
    .D(_00661_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _24129_ (.CLK(clknet_leaf_119_clk),
    .D(_00662_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[14] ));
 sky130_fd_sc_hd__dfxtp_2 _24130_ (.CLK(clknet_leaf_118_clk),
    .D(_00663_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[15] ));
 sky130_fd_sc_hd__dfxtp_2 _24131_ (.CLK(clknet_leaf_119_clk),
    .D(_00664_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[16] ));
 sky130_fd_sc_hd__dfxtp_1 _24132_ (.CLK(clknet_leaf_4_clk),
    .D(_00665_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[17] ));
 sky130_fd_sc_hd__dfxtp_1 _24133_ (.CLK(clknet_leaf_0_clk),
    .D(_00666_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[18] ));
 sky130_fd_sc_hd__dfxtp_1 _24134_ (.CLK(clknet_leaf_0_clk),
    .D(_00667_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[19] ));
 sky130_fd_sc_hd__dfxtp_1 _24135_ (.CLK(clknet_leaf_144_clk),
    .D(_00668_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[20] ));
 sky130_fd_sc_hd__dfxtp_1 _24136_ (.CLK(clknet_leaf_144_clk),
    .D(_00669_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[21] ));
 sky130_fd_sc_hd__dfxtp_1 _24137_ (.CLK(clknet_leaf_144_clk),
    .D(_00670_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[23] ));
 sky130_fd_sc_hd__dfxtp_1 _24138_ (.CLK(clknet_leaf_144_clk),
    .D(_00671_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[24] ));
 sky130_fd_sc_hd__dfxtp_2 _24139_ (.CLK(clknet_leaf_4_clk),
    .D(_00672_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[25] ));
 sky130_fd_sc_hd__dfxtp_1 _24140_ (.CLK(clknet_leaf_144_clk),
    .D(_00673_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[27] ));
 sky130_fd_sc_hd__dfxtp_1 _24141_ (.CLK(clknet_leaf_144_clk),
    .D(_00674_),
    .Q(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[31] ));
 sky130_fd_sc_hd__dfxtp_1 _24142_ (.CLK(clknet_leaf_14_clk),
    .D(_00675_),
    .Q(\top_inst.grid_inst.data_path_wires[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 _24143_ (.CLK(clknet_leaf_18_clk),
    .D(_00676_),
    .Q(\top_inst.grid_inst.data_path_wires[13][1] ));
 sky130_fd_sc_hd__dfxtp_2 _24144_ (.CLK(clknet_leaf_18_clk),
    .D(_00677_),
    .Q(\top_inst.grid_inst.data_path_wires[13][2] ));
 sky130_fd_sc_hd__dfxtp_2 _24145_ (.CLK(clknet_leaf_18_clk),
    .D(_00678_),
    .Q(\top_inst.grid_inst.data_path_wires[13][3] ));
 sky130_fd_sc_hd__dfxtp_2 _24146_ (.CLK(clknet_leaf_16_clk),
    .D(_00679_),
    .Q(\top_inst.grid_inst.data_path_wires[13][4] ));
 sky130_fd_sc_hd__dfxtp_2 _24147_ (.CLK(clknet_leaf_16_clk),
    .D(_00680_),
    .Q(\top_inst.grid_inst.data_path_wires[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 _24148_ (.CLK(clknet_leaf_16_clk),
    .D(_00681_),
    .Q(\top_inst.grid_inst.data_path_wires[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _24149_ (.CLK(clknet_leaf_17_clk),
    .D(_00682_),
    .Q(\top_inst.grid_inst.data_path_wires[13][7] ));
 sky130_fd_sc_hd__dfxtp_2 _24150_ (.CLK(clknet_leaf_18_clk),
    .D(_00683_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _24151_ (.CLK(clknet_leaf_18_clk),
    .D(_00684_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24152_ (.CLK(clknet_leaf_18_clk),
    .D(_00685_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _24153_ (.CLK(clknet_leaf_18_clk),
    .D(_00686_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _24154_ (.CLK(clknet_leaf_18_clk),
    .D(_00687_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24155_ (.CLK(clknet_leaf_18_clk),
    .D(_00688_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _24156_ (.CLK(clknet_leaf_17_clk),
    .D(_00689_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _24157_ (.CLK(clknet_leaf_17_clk),
    .D(_00690_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24158_ (.CLK(clknet_leaf_9_clk),
    .D(_00691_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[0] ));
 sky130_fd_sc_hd__dfxtp_1 _24159_ (.CLK(clknet_leaf_9_clk),
    .D(_00692_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24160_ (.CLK(clknet_leaf_9_clk),
    .D(_00693_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _24161_ (.CLK(clknet_leaf_13_clk),
    .D(_00694_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[3] ));
 sky130_fd_sc_hd__dfxtp_2 _24162_ (.CLK(clknet_leaf_13_clk),
    .D(_00695_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24163_ (.CLK(clknet_leaf_9_clk),
    .D(_00696_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[5] ));
 sky130_fd_sc_hd__dfxtp_1 _24164_ (.CLK(clknet_leaf_9_clk),
    .D(_00697_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[6] ));
 sky130_fd_sc_hd__dfxtp_2 _24165_ (.CLK(clknet_leaf_9_clk),
    .D(_00698_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[7] ));
 sky130_fd_sc_hd__dfxtp_2 _24166_ (.CLK(clknet_leaf_9_clk),
    .D(_00699_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[8] ));
 sky130_fd_sc_hd__dfxtp_1 _24167_ (.CLK(clknet_leaf_8_clk),
    .D(_00700_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[9] ));
 sky130_fd_sc_hd__dfxtp_2 _24168_ (.CLK(clknet_leaf_8_clk),
    .D(_00701_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[10] ));
 sky130_fd_sc_hd__dfxtp_1 _24169_ (.CLK(clknet_leaf_23_clk),
    .D(_00702_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[11] ));
 sky130_fd_sc_hd__dfxtp_1 _24170_ (.CLK(clknet_leaf_23_clk),
    .D(_00703_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[12] ));
 sky130_fd_sc_hd__dfxtp_1 _24171_ (.CLK(clknet_leaf_23_clk),
    .D(_00704_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _24172_ (.CLK(clknet_leaf_23_clk),
    .D(_00705_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[14] ));
 sky130_fd_sc_hd__dfxtp_1 _24173_ (.CLK(clknet_leaf_23_clk),
    .D(_00706_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[15] ));
 sky130_fd_sc_hd__dfxtp_1 _24174_ (.CLK(clknet_leaf_23_clk),
    .D(_00707_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[16] ));
 sky130_fd_sc_hd__dfxtp_1 _24175_ (.CLK(clknet_leaf_27_clk),
    .D(_00708_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[17] ));
 sky130_fd_sc_hd__dfxtp_1 _24176_ (.CLK(clknet_leaf_27_clk),
    .D(_00709_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[18] ));
 sky130_fd_sc_hd__dfxtp_1 _24177_ (.CLK(clknet_leaf_29_clk),
    .D(_00710_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[19] ));
 sky130_fd_sc_hd__dfxtp_1 _24178_ (.CLK(clknet_leaf_29_clk),
    .D(_00711_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[20] ));
 sky130_fd_sc_hd__dfxtp_1 _24179_ (.CLK(clknet_leaf_29_clk),
    .D(_00712_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[21] ));
 sky130_fd_sc_hd__dfxtp_1 _24180_ (.CLK(clknet_leaf_29_clk),
    .D(_00713_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[23] ));
 sky130_fd_sc_hd__dfxtp_1 _24181_ (.CLK(clknet_leaf_29_clk),
    .D(_00714_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[24] ));
 sky130_fd_sc_hd__dfxtp_2 _24182_ (.CLK(clknet_leaf_29_clk),
    .D(_00715_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[25] ));
 sky130_fd_sc_hd__dfxtp_1 _24183_ (.CLK(clknet_leaf_29_clk),
    .D(_00716_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[27] ));
 sky130_fd_sc_hd__dfxtp_1 _24184_ (.CLK(clknet_leaf_29_clk),
    .D(_00717_),
    .Q(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[31] ));
 sky130_fd_sc_hd__dfxtp_1 _24185_ (.CLK(clknet_leaf_47_clk),
    .D(_00718_),
    .Q(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _24186_ (.CLK(clknet_leaf_47_clk),
    .D(_00719_),
    .Q(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _24187_ (.CLK(clknet_leaf_47_clk),
    .D(_00720_),
    .Q(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _24188_ (.CLK(clknet_leaf_47_clk),
    .D(_00721_),
    .Q(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _24189_ (.CLK(clknet_leaf_47_clk),
    .D(_00722_),
    .Q(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24190_ (.CLK(clknet_leaf_48_clk),
    .D(_00723_),
    .Q(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _24191_ (.CLK(clknet_leaf_47_clk),
    .D(_00724_),
    .Q(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24192_ (.CLK(clknet_leaf_47_clk),
    .D(_00725_),
    .Q(\top_inst.grid_inst.rows[3].cols[0].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24193_ (.CLK(clknet_leaf_117_clk),
    .D(_00726_),
    .Q(\top_inst.deskew_buff_inst.col_input[0] ));
 sky130_fd_sc_hd__dfxtp_1 _24194_ (.CLK(clknet_leaf_117_clk),
    .D(_00727_),
    .Q(\top_inst.deskew_buff_inst.col_input[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24195_ (.CLK(clknet_leaf_15_clk),
    .D(_00728_),
    .Q(\top_inst.deskew_buff_inst.col_input[2] ));
 sky130_fd_sc_hd__dfxtp_1 _24196_ (.CLK(clknet_leaf_15_clk),
    .D(_00729_),
    .Q(\top_inst.deskew_buff_inst.col_input[3] ));
 sky130_fd_sc_hd__dfxtp_1 _24197_ (.CLK(clknet_leaf_15_clk),
    .D(_00730_),
    .Q(\top_inst.deskew_buff_inst.col_input[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24198_ (.CLK(clknet_leaf_116_clk),
    .D(_00731_),
    .Q(\top_inst.deskew_buff_inst.col_input[5] ));
 sky130_fd_sc_hd__dfxtp_1 _24199_ (.CLK(clknet_leaf_116_clk),
    .D(_00732_),
    .Q(\top_inst.deskew_buff_inst.col_input[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24200_ (.CLK(clknet_leaf_117_clk),
    .D(_00733_),
    .Q(\top_inst.deskew_buff_inst.col_input[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24201_ (.CLK(clknet_leaf_116_clk),
    .D(_00734_),
    .Q(\top_inst.deskew_buff_inst.col_input[8] ));
 sky130_fd_sc_hd__dfxtp_1 _24202_ (.CLK(clknet_leaf_117_clk),
    .D(_00735_),
    .Q(\top_inst.deskew_buff_inst.col_input[9] ));
 sky130_fd_sc_hd__dfxtp_1 _24203_ (.CLK(clknet_leaf_16_clk),
    .D(_00736_),
    .Q(\top_inst.deskew_buff_inst.col_input[10] ));
 sky130_fd_sc_hd__dfxtp_1 _24204_ (.CLK(clknet_leaf_16_clk),
    .D(_00737_),
    .Q(\top_inst.deskew_buff_inst.col_input[11] ));
 sky130_fd_sc_hd__dfxtp_1 _24205_ (.CLK(clknet_leaf_117_clk),
    .D(_00738_),
    .Q(\top_inst.deskew_buff_inst.col_input[12] ));
 sky130_fd_sc_hd__dfxtp_1 _24206_ (.CLK(clknet_leaf_117_clk),
    .D(_00739_),
    .Q(\top_inst.deskew_buff_inst.col_input[13] ));
 sky130_fd_sc_hd__dfxtp_1 _24207_ (.CLK(clknet_leaf_17_clk),
    .D(_00740_),
    .Q(\top_inst.deskew_buff_inst.col_input[14] ));
 sky130_fd_sc_hd__dfxtp_1 _24208_ (.CLK(clknet_leaf_17_clk),
    .D(_00741_),
    .Q(\top_inst.deskew_buff_inst.col_input[15] ));
 sky130_fd_sc_hd__dfxtp_1 _24209_ (.CLK(clknet_leaf_118_clk),
    .D(_00742_),
    .Q(\top_inst.deskew_buff_inst.col_input[16] ));
 sky130_fd_sc_hd__dfxtp_1 _24210_ (.CLK(clknet_leaf_17_clk),
    .D(_00743_),
    .Q(\top_inst.deskew_buff_inst.col_input[17] ));
 sky130_fd_sc_hd__dfxtp_1 _24211_ (.CLK(clknet_leaf_17_clk),
    .D(_00744_),
    .Q(\top_inst.deskew_buff_inst.col_input[18] ));
 sky130_fd_sc_hd__dfxtp_1 _24212_ (.CLK(clknet_leaf_118_clk),
    .D(_00745_),
    .Q(\top_inst.deskew_buff_inst.col_input[19] ));
 sky130_fd_sc_hd__dfxtp_1 _24213_ (.CLK(clknet_leaf_118_clk),
    .D(_00746_),
    .Q(\top_inst.deskew_buff_inst.col_input[20] ));
 sky130_fd_sc_hd__dfxtp_1 _24214_ (.CLK(clknet_leaf_17_clk),
    .D(_00747_),
    .Q(\top_inst.deskew_buff_inst.col_input[21] ));
 sky130_fd_sc_hd__dfxtp_1 _24215_ (.CLK(clknet_leaf_118_clk),
    .D(_00748_),
    .Q(\top_inst.deskew_buff_inst.col_input[22] ));
 sky130_fd_sc_hd__dfxtp_1 _24216_ (.CLK(clknet_leaf_19_clk),
    .D(_00749_),
    .Q(\top_inst.deskew_buff_inst.col_input[23] ));
 sky130_fd_sc_hd__dfxtp_1 _24217_ (.CLK(clknet_leaf_118_clk),
    .D(_00750_),
    .Q(\top_inst.deskew_buff_inst.col_input[24] ));
 sky130_fd_sc_hd__dfxtp_1 _24218_ (.CLK(clknet_leaf_19_clk),
    .D(_00751_),
    .Q(\top_inst.deskew_buff_inst.col_input[25] ));
 sky130_fd_sc_hd__dfxtp_1 _24219_ (.CLK(clknet_leaf_19_clk),
    .D(_00752_),
    .Q(\top_inst.deskew_buff_inst.col_input[26] ));
 sky130_fd_sc_hd__dfxtp_1 _24220_ (.CLK(clknet_leaf_19_clk),
    .D(_00753_),
    .Q(\top_inst.deskew_buff_inst.col_input[27] ));
 sky130_fd_sc_hd__dfxtp_1 _24221_ (.CLK(clknet_leaf_118_clk),
    .D(_00754_),
    .Q(\top_inst.deskew_buff_inst.col_input[28] ));
 sky130_fd_sc_hd__dfxtp_1 _24222_ (.CLK(clknet_leaf_12_clk),
    .D(_00755_),
    .Q(\top_inst.deskew_buff_inst.col_input[29] ));
 sky130_fd_sc_hd__dfxtp_1 _24223_ (.CLK(clknet_leaf_19_clk),
    .D(_00756_),
    .Q(\top_inst.deskew_buff_inst.col_input[30] ));
 sky130_fd_sc_hd__dfxtp_1 _24224_ (.CLK(clknet_leaf_19_clk),
    .D(_00757_),
    .Q(\top_inst.deskew_buff_inst.col_input[31] ));
 sky130_fd_sc_hd__dfxtp_1 _24225_ (.CLK(clknet_leaf_112_clk),
    .D(_00758_),
    .Q(\top_inst.grid_inst.data_path_wires[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _24226_ (.CLK(clknet_leaf_112_clk),
    .D(_00759_),
    .Q(\top_inst.grid_inst.data_path_wires[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _24227_ (.CLK(clknet_leaf_113_clk),
    .D(_00760_),
    .Q(\top_inst.grid_inst.data_path_wires[16][2] ));
 sky130_fd_sc_hd__dfxtp_2 _24228_ (.CLK(clknet_leaf_112_clk),
    .D(_00761_),
    .Q(\top_inst.grid_inst.data_path_wires[16][3] ));
 sky130_fd_sc_hd__dfxtp_4 _24229_ (.CLK(clknet_leaf_113_clk),
    .D(_00762_),
    .Q(\top_inst.grid_inst.data_path_wires[16][4] ));
 sky130_fd_sc_hd__dfxtp_2 _24230_ (.CLK(clknet_leaf_113_clk),
    .D(_00763_),
    .Q(\top_inst.grid_inst.data_path_wires[16][5] ));
 sky130_fd_sc_hd__dfxtp_4 _24231_ (.CLK(clknet_leaf_113_clk),
    .D(_00764_),
    .Q(\top_inst.grid_inst.data_path_wires[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _24232_ (.CLK(clknet_leaf_111_clk),
    .D(_00765_),
    .Q(\top_inst.grid_inst.data_path_wires[16][7] ));
 sky130_fd_sc_hd__dfxtp_2 _24233_ (.CLK(clknet_leaf_112_clk),
    .D(_00766_),
    .Q(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _24234_ (.CLK(clknet_leaf_112_clk),
    .D(_00767_),
    .Q(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24235_ (.CLK(clknet_leaf_113_clk),
    .D(_00768_),
    .Q(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_4 _24236_ (.CLK(clknet_leaf_113_clk),
    .D(_00769_),
    .Q(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _24237_ (.CLK(clknet_leaf_113_clk),
    .D(_00770_),
    .Q(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24238_ (.CLK(clknet_leaf_111_clk),
    .D(_00771_),
    .Q(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _24239_ (.CLK(clknet_leaf_111_clk),
    .D(_00772_),
    .Q(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _24240_ (.CLK(clknet_leaf_113_clk),
    .D(_00773_),
    .Q(\top_inst.grid_inst.rows[3].cols[1].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24241_ (.CLK(clknet_leaf_112_clk),
    .D(_00774_),
    .Q(\top_inst.deskew_buff_inst.col_input[32] ));
 sky130_fd_sc_hd__dfxtp_1 _24242_ (.CLK(clknet_leaf_108_clk),
    .D(_00775_),
    .Q(\top_inst.deskew_buff_inst.col_input[33] ));
 sky130_fd_sc_hd__dfxtp_1 _24243_ (.CLK(clknet_leaf_116_clk),
    .D(_00776_),
    .Q(\top_inst.deskew_buff_inst.col_input[34] ));
 sky130_fd_sc_hd__dfxtp_1 _24244_ (.CLK(clknet_leaf_125_clk),
    .D(_00777_),
    .Q(\top_inst.deskew_buff_inst.col_input[35] ));
 sky130_fd_sc_hd__dfxtp_1 _24245_ (.CLK(clknet_leaf_126_clk),
    .D(_00778_),
    .Q(\top_inst.deskew_buff_inst.col_input[36] ));
 sky130_fd_sc_hd__dfxtp_1 _24246_ (.CLK(clknet_leaf_108_clk),
    .D(_00779_),
    .Q(\top_inst.deskew_buff_inst.col_input[37] ));
 sky130_fd_sc_hd__dfxtp_1 _24247_ (.CLK(clknet_leaf_108_clk),
    .D(_00780_),
    .Q(\top_inst.deskew_buff_inst.col_input[38] ));
 sky130_fd_sc_hd__dfxtp_1 _24248_ (.CLK(clknet_leaf_108_clk),
    .D(_00781_),
    .Q(\top_inst.deskew_buff_inst.col_input[39] ));
 sky130_fd_sc_hd__dfxtp_1 _24249_ (.CLK(clknet_leaf_107_clk),
    .D(_00782_),
    .Q(\top_inst.deskew_buff_inst.col_input[40] ));
 sky130_fd_sc_hd__dfxtp_1 _24250_ (.CLK(clknet_leaf_108_clk),
    .D(_00783_),
    .Q(\top_inst.deskew_buff_inst.col_input[41] ));
 sky130_fd_sc_hd__dfxtp_1 _24251_ (.CLK(clknet_leaf_107_clk),
    .D(_00784_),
    .Q(\top_inst.deskew_buff_inst.col_input[42] ));
 sky130_fd_sc_hd__dfxtp_1 _24252_ (.CLK(clknet_leaf_107_clk),
    .D(_00785_),
    .Q(\top_inst.deskew_buff_inst.col_input[43] ));
 sky130_fd_sc_hd__dfxtp_1 _24253_ (.CLK(clknet_leaf_106_clk),
    .D(_00786_),
    .Q(\top_inst.deskew_buff_inst.col_input[44] ));
 sky130_fd_sc_hd__dfxtp_1 _24254_ (.CLK(clknet_leaf_110_clk),
    .D(_00787_),
    .Q(\top_inst.deskew_buff_inst.col_input[45] ));
 sky130_fd_sc_hd__dfxtp_1 _24255_ (.CLK(clknet_leaf_110_clk),
    .D(_00788_),
    .Q(\top_inst.deskew_buff_inst.col_input[46] ));
 sky130_fd_sc_hd__dfxtp_1 _24256_ (.CLK(clknet_leaf_110_clk),
    .D(_00789_),
    .Q(\top_inst.deskew_buff_inst.col_input[47] ));
 sky130_fd_sc_hd__dfxtp_1 _24257_ (.CLK(clknet_leaf_110_clk),
    .D(_00790_),
    .Q(\top_inst.deskew_buff_inst.col_input[48] ));
 sky130_fd_sc_hd__dfxtp_1 _24258_ (.CLK(clknet_leaf_110_clk),
    .D(_00791_),
    .Q(\top_inst.deskew_buff_inst.col_input[49] ));
 sky130_fd_sc_hd__dfxtp_1 _24259_ (.CLK(clknet_leaf_110_clk),
    .D(_00792_),
    .Q(\top_inst.deskew_buff_inst.col_input[50] ));
 sky130_fd_sc_hd__dfxtp_1 _24260_ (.CLK(clknet_leaf_110_clk),
    .D(_00793_),
    .Q(\top_inst.deskew_buff_inst.col_input[51] ));
 sky130_fd_sc_hd__dfxtp_1 _24261_ (.CLK(clknet_leaf_110_clk),
    .D(_00794_),
    .Q(\top_inst.deskew_buff_inst.col_input[52] ));
 sky130_fd_sc_hd__dfxtp_1 _24262_ (.CLK(clknet_leaf_110_clk),
    .D(_00795_),
    .Q(\top_inst.deskew_buff_inst.col_input[53] ));
 sky130_fd_sc_hd__dfxtp_1 _24263_ (.CLK(clknet_leaf_110_clk),
    .D(_00796_),
    .Q(\top_inst.deskew_buff_inst.col_input[54] ));
 sky130_fd_sc_hd__dfxtp_1 _24264_ (.CLK(clknet_leaf_105_clk),
    .D(_00797_),
    .Q(\top_inst.deskew_buff_inst.col_input[55] ));
 sky130_fd_sc_hd__dfxtp_1 _24265_ (.CLK(clknet_leaf_101_clk),
    .D(_00798_),
    .Q(\top_inst.deskew_buff_inst.col_input[56] ));
 sky130_fd_sc_hd__dfxtp_1 _24266_ (.CLK(clknet_leaf_100_clk),
    .D(_00799_),
    .Q(\top_inst.deskew_buff_inst.col_input[57] ));
 sky130_fd_sc_hd__dfxtp_1 _24267_ (.CLK(clknet_leaf_101_clk),
    .D(_00800_),
    .Q(\top_inst.deskew_buff_inst.col_input[58] ));
 sky130_fd_sc_hd__dfxtp_1 _24268_ (.CLK(clknet_leaf_100_clk),
    .D(_00801_),
    .Q(\top_inst.deskew_buff_inst.col_input[59] ));
 sky130_fd_sc_hd__dfxtp_1 _24269_ (.CLK(clknet_leaf_105_clk),
    .D(_00802_),
    .Q(\top_inst.deskew_buff_inst.col_input[60] ));
 sky130_fd_sc_hd__dfxtp_1 _24270_ (.CLK(clknet_leaf_100_clk),
    .D(_00803_),
    .Q(\top_inst.deskew_buff_inst.col_input[61] ));
 sky130_fd_sc_hd__dfxtp_1 _24271_ (.CLK(clknet_leaf_97_clk),
    .D(_00804_),
    .Q(\top_inst.deskew_buff_inst.col_input[62] ));
 sky130_fd_sc_hd__dfxtp_1 _24272_ (.CLK(clknet_leaf_97_clk),
    .D(_00805_),
    .Q(\top_inst.deskew_buff_inst.col_input[63] ));
 sky130_fd_sc_hd__dfxtp_1 _24273_ (.CLK(clknet_leaf_11_clk),
    .D(_00806_),
    .Q(\top_inst.grid_inst.data_path_wires[17][0] ));
 sky130_fd_sc_hd__dfxtp_2 _24274_ (.CLK(clknet_leaf_12_clk),
    .D(_00807_),
    .Q(\top_inst.grid_inst.data_path_wires[17][1] ));
 sky130_fd_sc_hd__dfxtp_2 _24275_ (.CLK(clknet_leaf_11_clk),
    .D(_00808_),
    .Q(\top_inst.grid_inst.data_path_wires[17][2] ));
 sky130_fd_sc_hd__dfxtp_2 _24276_ (.CLK(clknet_leaf_11_clk),
    .D(_00809_),
    .Q(\top_inst.grid_inst.data_path_wires[17][3] ));
 sky130_fd_sc_hd__dfxtp_2 _24277_ (.CLK(clknet_leaf_11_clk),
    .D(_00810_),
    .Q(\top_inst.grid_inst.data_path_wires[17][4] ));
 sky130_fd_sc_hd__dfxtp_2 _24278_ (.CLK(clknet_leaf_12_clk),
    .D(_00811_),
    .Q(\top_inst.grid_inst.data_path_wires[17][5] ));
 sky130_fd_sc_hd__dfxtp_2 _24279_ (.CLK(clknet_leaf_11_clk),
    .D(_00812_),
    .Q(\top_inst.grid_inst.data_path_wires[17][6] ));
 sky130_fd_sc_hd__dfxtp_2 _24280_ (.CLK(clknet_leaf_11_clk),
    .D(_00813_),
    .Q(\top_inst.grid_inst.data_path_wires[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _24281_ (.CLK(clknet_leaf_11_clk),
    .D(_00814_),
    .Q(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _24282_ (.CLK(clknet_leaf_13_clk),
    .D(_00815_),
    .Q(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _24283_ (.CLK(clknet_leaf_10_clk),
    .D(_00816_),
    .Q(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _24284_ (.CLK(clknet_leaf_10_clk),
    .D(_00817_),
    .Q(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _24285_ (.CLK(clknet_leaf_10_clk),
    .D(_00818_),
    .Q(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24286_ (.CLK(clknet_4_4__leaf_clk),
    .D(_00819_),
    .Q(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _24287_ (.CLK(clknet_leaf_10_clk),
    .D(_00820_),
    .Q(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24288_ (.CLK(clknet_leaf_10_clk),
    .D(_00821_),
    .Q(\top_inst.grid_inst.rows[3].cols[2].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24289_ (.CLK(clknet_leaf_12_clk),
    .D(_00822_),
    .Q(\top_inst.deskew_buff_inst.col_input[64] ));
 sky130_fd_sc_hd__dfxtp_1 _24290_ (.CLK(clknet_leaf_120_clk),
    .D(_00823_),
    .Q(\top_inst.deskew_buff_inst.col_input[65] ));
 sky130_fd_sc_hd__dfxtp_1 _24291_ (.CLK(clknet_leaf_120_clk),
    .D(_00824_),
    .Q(\top_inst.deskew_buff_inst.col_input[66] ));
 sky130_fd_sc_hd__dfxtp_1 _24292_ (.CLK(clknet_leaf_120_clk),
    .D(_00825_),
    .Q(\top_inst.deskew_buff_inst.col_input[67] ));
 sky130_fd_sc_hd__dfxtp_1 _24293_ (.CLK(clknet_leaf_120_clk),
    .D(_00826_),
    .Q(\top_inst.deskew_buff_inst.col_input[68] ));
 sky130_fd_sc_hd__dfxtp_1 _24294_ (.CLK(clknet_leaf_137_clk),
    .D(_00827_),
    .Q(\top_inst.deskew_buff_inst.col_input[69] ));
 sky130_fd_sc_hd__dfxtp_1 _24295_ (.CLK(clknet_leaf_137_clk),
    .D(_00828_),
    .Q(\top_inst.deskew_buff_inst.col_input[70] ));
 sky130_fd_sc_hd__dfxtp_1 _24296_ (.CLK(clknet_leaf_137_clk),
    .D(_00829_),
    .Q(\top_inst.deskew_buff_inst.col_input[71] ));
 sky130_fd_sc_hd__dfxtp_1 _24297_ (.CLK(clknet_leaf_137_clk),
    .D(_00830_),
    .Q(\top_inst.deskew_buff_inst.col_input[72] ));
 sky130_fd_sc_hd__dfxtp_1 _24298_ (.CLK(clknet_leaf_137_clk),
    .D(_00831_),
    .Q(\top_inst.deskew_buff_inst.col_input[73] ));
 sky130_fd_sc_hd__dfxtp_1 _24299_ (.CLK(clknet_leaf_138_clk),
    .D(_00832_),
    .Q(\top_inst.deskew_buff_inst.col_input[74] ));
 sky130_fd_sc_hd__dfxtp_1 _24300_ (.CLK(clknet_leaf_138_clk),
    .D(_00833_),
    .Q(\top_inst.deskew_buff_inst.col_input[75] ));
 sky130_fd_sc_hd__dfxtp_1 _24301_ (.CLK(clknet_leaf_138_clk),
    .D(_00834_),
    .Q(\top_inst.deskew_buff_inst.col_input[76] ));
 sky130_fd_sc_hd__dfxtp_1 _24302_ (.CLK(clknet_leaf_138_clk),
    .D(_00835_),
    .Q(\top_inst.deskew_buff_inst.col_input[77] ));
 sky130_fd_sc_hd__dfxtp_1 _24303_ (.CLK(clknet_leaf_2_clk),
    .D(_00836_),
    .Q(\top_inst.deskew_buff_inst.col_input[78] ));
 sky130_fd_sc_hd__dfxtp_1 _24304_ (.CLK(clknet_leaf_2_clk),
    .D(_00837_),
    .Q(\top_inst.deskew_buff_inst.col_input[79] ));
 sky130_fd_sc_hd__dfxtp_1 _24305_ (.CLK(clknet_leaf_2_clk),
    .D(_00838_),
    .Q(\top_inst.deskew_buff_inst.col_input[80] ));
 sky130_fd_sc_hd__dfxtp_1 _24306_ (.CLK(clknet_leaf_138_clk),
    .D(_00839_),
    .Q(\top_inst.deskew_buff_inst.col_input[81] ));
 sky130_fd_sc_hd__dfxtp_1 _24307_ (.CLK(clknet_leaf_2_clk),
    .D(_00840_),
    .Q(\top_inst.deskew_buff_inst.col_input[82] ));
 sky130_fd_sc_hd__dfxtp_1 _24308_ (.CLK(clknet_leaf_2_clk),
    .D(_00841_),
    .Q(\top_inst.deskew_buff_inst.col_input[83] ));
 sky130_fd_sc_hd__dfxtp_1 _24309_ (.CLK(clknet_leaf_1_clk),
    .D(_00842_),
    .Q(\top_inst.deskew_buff_inst.col_input[84] ));
 sky130_fd_sc_hd__dfxtp_1 _24310_ (.CLK(clknet_leaf_2_clk),
    .D(_00843_),
    .Q(\top_inst.deskew_buff_inst.col_input[85] ));
 sky130_fd_sc_hd__dfxtp_1 _24311_ (.CLK(clknet_leaf_2_clk),
    .D(_00844_),
    .Q(\top_inst.deskew_buff_inst.col_input[86] ));
 sky130_fd_sc_hd__dfxtp_1 _24312_ (.CLK(clknet_leaf_1_clk),
    .D(_00845_),
    .Q(\top_inst.deskew_buff_inst.col_input[87] ));
 sky130_fd_sc_hd__dfxtp_1 _24313_ (.CLK(clknet_leaf_1_clk),
    .D(_00846_),
    .Q(\top_inst.deskew_buff_inst.col_input[88] ));
 sky130_fd_sc_hd__dfxtp_1 _24314_ (.CLK(clknet_leaf_1_clk),
    .D(_00847_),
    .Q(\top_inst.deskew_buff_inst.col_input[89] ));
 sky130_fd_sc_hd__dfxtp_1 _24315_ (.CLK(clknet_leaf_1_clk),
    .D(_00848_),
    .Q(\top_inst.deskew_buff_inst.col_input[90] ));
 sky130_fd_sc_hd__dfxtp_1 _24316_ (.CLK(clknet_leaf_1_clk),
    .D(_00849_),
    .Q(\top_inst.deskew_buff_inst.col_input[91] ));
 sky130_fd_sc_hd__dfxtp_1 _24317_ (.CLK(clknet_leaf_1_clk),
    .D(_00850_),
    .Q(\top_inst.deskew_buff_inst.col_input[92] ));
 sky130_fd_sc_hd__dfxtp_1 _24318_ (.CLK(clknet_leaf_2_clk),
    .D(_00851_),
    .Q(\top_inst.deskew_buff_inst.col_input[93] ));
 sky130_fd_sc_hd__dfxtp_1 _24319_ (.CLK(clknet_leaf_139_clk),
    .D(_00852_),
    .Q(\top_inst.deskew_buff_inst.col_input[94] ));
 sky130_fd_sc_hd__dfxtp_1 _24320_ (.CLK(clknet_leaf_143_clk),
    .D(_00853_),
    .Q(\top_inst.deskew_buff_inst.col_input[95] ));
 sky130_fd_sc_hd__dfxtp_2 _24321_ (.CLK(clknet_leaf_9_clk),
    .D(_00854_),
    .Q(\top_inst.grid_inst.data_path_wires[18][0] ));
 sky130_fd_sc_hd__dfxtp_2 _24322_ (.CLK(clknet_leaf_10_clk),
    .D(_00855_),
    .Q(\top_inst.grid_inst.data_path_wires[18][1] ));
 sky130_fd_sc_hd__dfxtp_2 _24323_ (.CLK(clknet_leaf_5_clk),
    .D(_00856_),
    .Q(\top_inst.grid_inst.data_path_wires[18][2] ));
 sky130_fd_sc_hd__dfxtp_2 _24324_ (.CLK(clknet_leaf_10_clk),
    .D(_00857_),
    .Q(\top_inst.grid_inst.data_path_wires[18][3] ));
 sky130_fd_sc_hd__dfxtp_2 _24325_ (.CLK(clknet_leaf_10_clk),
    .D(_00858_),
    .Q(\top_inst.grid_inst.data_path_wires[18][4] ));
 sky130_fd_sc_hd__dfxtp_2 _24326_ (.CLK(clknet_leaf_7_clk),
    .D(_00859_),
    .Q(\top_inst.grid_inst.data_path_wires[18][5] ));
 sky130_fd_sc_hd__dfxtp_2 _24327_ (.CLK(clknet_leaf_5_clk),
    .D(_00860_),
    .Q(\top_inst.grid_inst.data_path_wires[18][6] ));
 sky130_fd_sc_hd__dfxtp_4 _24328_ (.CLK(clknet_leaf_5_clk),
    .D(_00861_),
    .Q(\top_inst.grid_inst.data_path_wires[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _24329_ (.CLK(clknet_leaf_6_clk),
    .D(_00862_),
    .Q(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _24330_ (.CLK(clknet_leaf_7_clk),
    .D(_00863_),
    .Q(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24331_ (.CLK(clknet_leaf_6_clk),
    .D(_00864_),
    .Q(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _24332_ (.CLK(clknet_leaf_5_clk),
    .D(_00865_),
    .Q(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _24333_ (.CLK(clknet_leaf_5_clk),
    .D(_00866_),
    .Q(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _24334_ (.CLK(clknet_leaf_5_clk),
    .D(_00867_),
    .Q(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _24335_ (.CLK(clknet_leaf_5_clk),
    .D(_00868_),
    .Q(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24336_ (.CLK(clknet_leaf_5_clk),
    .D(_00869_),
    .Q(\top_inst.grid_inst.rows[3].cols[3].pe_inst.weight_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24337_ (.CLK(clknet_leaf_9_clk),
    .D(_00870_),
    .Q(\top_inst.deskew_buff_inst.col_input[96] ));
 sky130_fd_sc_hd__dfxtp_1 _24338_ (.CLK(clknet_leaf_9_clk),
    .D(_00871_),
    .Q(\top_inst.deskew_buff_inst.col_input[97] ));
 sky130_fd_sc_hd__dfxtp_1 _24339_ (.CLK(clknet_leaf_9_clk),
    .D(_00872_),
    .Q(\top_inst.deskew_buff_inst.col_input[98] ));
 sky130_fd_sc_hd__dfxtp_1 _24340_ (.CLK(clknet_leaf_8_clk),
    .D(_00873_),
    .Q(\top_inst.deskew_buff_inst.col_input[99] ));
 sky130_fd_sc_hd__dfxtp_1 _24341_ (.CLK(clknet_leaf_8_clk),
    .D(_00874_),
    .Q(\top_inst.deskew_buff_inst.col_input[100] ));
 sky130_fd_sc_hd__dfxtp_1 _24342_ (.CLK(clknet_leaf_8_clk),
    .D(_00875_),
    .Q(\top_inst.deskew_buff_inst.col_input[101] ));
 sky130_fd_sc_hd__dfxtp_1 _24343_ (.CLK(clknet_leaf_8_clk),
    .D(_00876_),
    .Q(\top_inst.deskew_buff_inst.col_input[102] ));
 sky130_fd_sc_hd__dfxtp_1 _24344_ (.CLK(clknet_leaf_8_clk),
    .D(_00877_),
    .Q(\top_inst.deskew_buff_inst.col_input[103] ));
 sky130_fd_sc_hd__dfxtp_1 _24345_ (.CLK(clknet_leaf_24_clk),
    .D(_00878_),
    .Q(\top_inst.deskew_buff_inst.col_input[104] ));
 sky130_fd_sc_hd__dfxtp_1 _24346_ (.CLK(clknet_leaf_24_clk),
    .D(_00879_),
    .Q(\top_inst.deskew_buff_inst.col_input[105] ));
 sky130_fd_sc_hd__dfxtp_1 _24347_ (.CLK(clknet_leaf_26_clk),
    .D(_00880_),
    .Q(\top_inst.deskew_buff_inst.col_input[106] ));
 sky130_fd_sc_hd__dfxtp_1 _24348_ (.CLK(clknet_leaf_24_clk),
    .D(_00881_),
    .Q(\top_inst.deskew_buff_inst.col_input[107] ));
 sky130_fd_sc_hd__dfxtp_1 _24349_ (.CLK(clknet_leaf_23_clk),
    .D(_00882_),
    .Q(\top_inst.deskew_buff_inst.col_input[108] ));
 sky130_fd_sc_hd__dfxtp_1 _24350_ (.CLK(clknet_leaf_24_clk),
    .D(_00883_),
    .Q(\top_inst.deskew_buff_inst.col_input[109] ));
 sky130_fd_sc_hd__dfxtp_1 _24351_ (.CLK(clknet_leaf_26_clk),
    .D(_00884_),
    .Q(\top_inst.deskew_buff_inst.col_input[110] ));
 sky130_fd_sc_hd__dfxtp_1 _24352_ (.CLK(clknet_leaf_24_clk),
    .D(_00885_),
    .Q(\top_inst.deskew_buff_inst.col_input[111] ));
 sky130_fd_sc_hd__dfxtp_1 _24353_ (.CLK(clknet_leaf_26_clk),
    .D(_00886_),
    .Q(\top_inst.deskew_buff_inst.col_input[112] ));
 sky130_fd_sc_hd__dfxtp_1 _24354_ (.CLK(clknet_leaf_26_clk),
    .D(_00887_),
    .Q(\top_inst.deskew_buff_inst.col_input[113] ));
 sky130_fd_sc_hd__dfxtp_1 _24355_ (.CLK(clknet_leaf_21_clk),
    .D(_00888_),
    .Q(\top_inst.deskew_buff_inst.col_input[114] ));
 sky130_fd_sc_hd__dfxtp_1 _24356_ (.CLK(clknet_leaf_26_clk),
    .D(_00889_),
    .Q(\top_inst.deskew_buff_inst.col_input[115] ));
 sky130_fd_sc_hd__dfxtp_1 _24357_ (.CLK(clknet_leaf_22_clk),
    .D(_00890_),
    .Q(\top_inst.deskew_buff_inst.col_input[116] ));
 sky130_fd_sc_hd__dfxtp_1 _24358_ (.CLK(clknet_4_5__leaf_clk),
    .D(_00891_),
    .Q(\top_inst.deskew_buff_inst.col_input[117] ));
 sky130_fd_sc_hd__dfxtp_1 _24359_ (.CLK(clknet_leaf_30_clk),
    .D(_00892_),
    .Q(\top_inst.deskew_buff_inst.col_input[118] ));
 sky130_fd_sc_hd__dfxtp_1 _24360_ (.CLK(clknet_leaf_30_clk),
    .D(_00893_),
    .Q(\top_inst.deskew_buff_inst.col_input[119] ));
 sky130_fd_sc_hd__dfxtp_1 _24361_ (.CLK(clknet_leaf_30_clk),
    .D(_00894_),
    .Q(\top_inst.deskew_buff_inst.col_input[120] ));
 sky130_fd_sc_hd__dfxtp_1 _24362_ (.CLK(clknet_leaf_30_clk),
    .D(_00895_),
    .Q(\top_inst.deskew_buff_inst.col_input[121] ));
 sky130_fd_sc_hd__dfxtp_1 _24363_ (.CLK(clknet_leaf_30_clk),
    .D(_00896_),
    .Q(\top_inst.deskew_buff_inst.col_input[122] ));
 sky130_fd_sc_hd__dfxtp_1 _24364_ (.CLK(clknet_leaf_31_clk),
    .D(_00897_),
    .Q(\top_inst.deskew_buff_inst.col_input[123] ));
 sky130_fd_sc_hd__dfxtp_1 _24365_ (.CLK(clknet_leaf_31_clk),
    .D(_00898_),
    .Q(\top_inst.deskew_buff_inst.col_input[124] ));
 sky130_fd_sc_hd__dfxtp_1 _24366_ (.CLK(clknet_leaf_31_clk),
    .D(_00899_),
    .Q(\top_inst.deskew_buff_inst.col_input[125] ));
 sky130_fd_sc_hd__dfxtp_1 _24367_ (.CLK(clknet_leaf_31_clk),
    .D(_00900_),
    .Q(\top_inst.deskew_buff_inst.col_input[126] ));
 sky130_fd_sc_hd__dfxtp_1 _24368_ (.CLK(clknet_leaf_31_clk),
    .D(_00901_),
    .Q(\top_inst.deskew_buff_inst.col_input[127] ));
 sky130_fd_sc_hd__dfxtp_1 _24369_ (.CLK(clknet_leaf_37_clk),
    .D(net937),
    .Q(\top_inst.skew_buff_inst.row[3].output_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _24370_ (.CLK(clknet_leaf_40_clk),
    .D(net579),
    .Q(\top_inst.skew_buff_inst.row[3].output_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24371_ (.CLK(clknet_leaf_37_clk),
    .D(net656),
    .Q(\top_inst.skew_buff_inst.row[3].output_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _24372_ (.CLK(clknet_leaf_39_clk),
    .D(net407),
    .Q(\top_inst.skew_buff_inst.row[3].output_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _24373_ (.CLK(clknet_leaf_38_clk),
    .D(net899),
    .Q(\top_inst.skew_buff_inst.row[3].output_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24374_ (.CLK(clknet_leaf_40_clk),
    .D(net675),
    .Q(\top_inst.skew_buff_inst.row[3].output_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _24375_ (.CLK(clknet_leaf_39_clk),
    .D(net395),
    .Q(\top_inst.skew_buff_inst.row[3].output_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24376_ (.CLK(clknet_leaf_39_clk),
    .D(net851),
    .Q(\top_inst.skew_buff_inst.row[3].output_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24377_ (.CLK(clknet_leaf_38_clk),
    .D(_00910_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _24378_ (.CLK(clknet_leaf_38_clk),
    .D(_00911_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _24379_ (.CLK(clknet_leaf_37_clk),
    .D(_00912_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _24380_ (.CLK(clknet_leaf_39_clk),
    .D(_00913_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _24381_ (.CLK(clknet_leaf_38_clk),
    .D(_00914_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _24382_ (.CLK(clknet_leaf_38_clk),
    .D(_00915_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _24383_ (.CLK(clknet_leaf_39_clk),
    .D(_00916_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _24384_ (.CLK(clknet_leaf_39_clk),
    .D(_00917_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _24385_ (.CLK(clknet_leaf_38_clk),
    .D(net716),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _24386_ (.CLK(clknet_leaf_38_clk),
    .D(_00919_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _24387_ (.CLK(clknet_leaf_38_clk),
    .D(net388),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _24388_ (.CLK(clknet_leaf_39_clk),
    .D(_00921_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _24389_ (.CLK(clknet_leaf_38_clk),
    .D(_00922_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _24390_ (.CLK(clknet_leaf_38_clk),
    .D(_00923_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _24391_ (.CLK(clknet_leaf_38_clk),
    .D(net295),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _24392_ (.CLK(clknet_leaf_39_clk),
    .D(net709),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _24393_ (.CLK(clknet_leaf_38_clk),
    .D(net853),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _24394_ (.CLK(clknet_leaf_38_clk),
    .D(_00927_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _24395_ (.CLK(clknet_leaf_37_clk),
    .D(_00928_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _24396_ (.CLK(clknet_leaf_38_clk),
    .D(net297),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _24397_ (.CLK(clknet_leaf_38_clk),
    .D(net785),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _24398_ (.CLK(clknet_leaf_38_clk),
    .D(_00931_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _24399_ (.CLK(clknet_leaf_38_clk),
    .D(_00932_),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _24400_ (.CLK(clknet_leaf_39_clk),
    .D(net765),
    .Q(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _24401_ (.CLK(clknet_leaf_57_clk),
    .D(net397),
    .Q(\top_inst.skew_buff_inst.row[2].output_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _24402_ (.CLK(clknet_leaf_57_clk),
    .D(net770),
    .Q(\top_inst.skew_buff_inst.row[2].output_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24403_ (.CLK(clknet_leaf_55_clk),
    .D(net767),
    .Q(\top_inst.skew_buff_inst.row[2].output_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _24404_ (.CLK(clknet_leaf_57_clk),
    .D(net414),
    .Q(\top_inst.skew_buff_inst.row[2].output_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _24405_ (.CLK(clknet_leaf_39_clk),
    .D(net417),
    .Q(\top_inst.skew_buff_inst.row[2].output_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24406_ (.CLK(clknet_leaf_57_clk),
    .D(net390),
    .Q(\top_inst.skew_buff_inst.row[2].output_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _24407_ (.CLK(clknet_leaf_55_clk),
    .D(net381),
    .Q(\top_inst.skew_buff_inst.row[2].output_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24408_ (.CLK(clknet_leaf_39_clk),
    .D(net713),
    .Q(\top_inst.skew_buff_inst.row[2].output_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24409_ (.CLK(clknet_leaf_57_clk),
    .D(_00942_),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _24410_ (.CLK(clknet_leaf_57_clk),
    .D(_00943_),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _24411_ (.CLK(clknet_leaf_55_clk),
    .D(_00944_),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _24412_ (.CLK(clknet_leaf_55_clk),
    .D(_00945_),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _24413_ (.CLK(clknet_leaf_56_clk),
    .D(net591),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _24414_ (.CLK(clknet_leaf_56_clk),
    .D(_00947_),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _24415_ (.CLK(clknet_leaf_56_clk),
    .D(_00948_),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _24416_ (.CLK(clknet_leaf_56_clk),
    .D(_00949_),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _24417_ (.CLK(clknet_leaf_56_clk),
    .D(_00950_),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _24418_ (.CLK(clknet_leaf_57_clk),
    .D(net644),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _24419_ (.CLK(clknet_leaf_55_clk),
    .D(net663),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _24420_ (.CLK(clknet_leaf_58_clk),
    .D(_00953_),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _24421_ (.CLK(clknet_leaf_56_clk),
    .D(_00954_),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _24422_ (.CLK(clknet_leaf_56_clk),
    .D(_00955_),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _24423_ (.CLK(clknet_leaf_56_clk),
    .D(_00956_),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _24424_ (.CLK(clknet_leaf_39_clk),
    .D(net405),
    .Q(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _24425_ (.CLK(clknet_leaf_57_clk),
    .D(net735),
    .Q(\top_inst.skew_buff_inst.row[1].output_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _24426_ (.CLK(clknet_leaf_58_clk),
    .D(net603),
    .Q(\top_inst.skew_buff_inst.row[1].output_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24427_ (.CLK(clknet_leaf_54_clk),
    .D(net773),
    .Q(\top_inst.skew_buff_inst.row[1].output_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _24428_ (.CLK(clknet_leaf_54_clk),
    .D(net703),
    .Q(\top_inst.skew_buff_inst.row[1].output_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _24429_ (.CLK(clknet_leaf_58_clk),
    .D(net719),
    .Q(\top_inst.skew_buff_inst.row[1].output_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24430_ (.CLK(clknet_leaf_59_clk),
    .D(net882),
    .Q(\top_inst.skew_buff_inst.row[1].output_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _24431_ (.CLK(clknet_leaf_58_clk),
    .D(net638),
    .Q(\top_inst.skew_buff_inst.row[1].output_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24432_ (.CLK(clknet_leaf_58_clk),
    .D(net634),
    .Q(\top_inst.skew_buff_inst.row[1].output_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24433_ (.CLK(clknet_leaf_57_clk),
    .D(net607),
    .Q(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _24434_ (.CLK(clknet_leaf_58_clk),
    .D(_00967_),
    .Q(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _24435_ (.CLK(clknet_leaf_54_clk),
    .D(_00968_),
    .Q(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _24436_ (.CLK(clknet_leaf_54_clk),
    .D(_00969_),
    .Q(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _24437_ (.CLK(clknet_leaf_58_clk),
    .D(_00970_),
    .Q(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _24438_ (.CLK(clknet_leaf_57_clk),
    .D(_00971_),
    .Q(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _24439_ (.CLK(clknet_leaf_58_clk),
    .D(net584),
    .Q(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _24440_ (.CLK(clknet_leaf_54_clk),
    .D(_00973_),
    .Q(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _24441_ (.CLK(clknet_leaf_64_clk),
    .D(net904),
    .Q(\top_inst.skew_buff_inst.row[0].output_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _24442_ (.CLK(clknet_leaf_64_clk),
    .D(net984),
    .Q(\top_inst.skew_buff_inst.row[0].output_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24443_ (.CLK(clknet_leaf_63_clk),
    .D(net952),
    .Q(\top_inst.skew_buff_inst.row[0].output_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _24444_ (.CLK(clknet_leaf_64_clk),
    .D(net980),
    .Q(\top_inst.skew_buff_inst.row[0].output_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _24445_ (.CLK(clknet_leaf_63_clk),
    .D(net1020),
    .Q(\top_inst.skew_buff_inst.row[0].output_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24446_ (.CLK(clknet_leaf_63_clk),
    .D(net617),
    .Q(\top_inst.skew_buff_inst.row[0].output_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _24447_ (.CLK(clknet_leaf_63_clk),
    .D(_00980_),
    .Q(\top_inst.skew_buff_inst.row[0].output_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24448_ (.CLK(clknet_leaf_63_clk),
    .D(net259),
    .Q(\top_inst.skew_buff_inst.row[0].output_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24449_ (.CLK(clknet_leaf_63_clk),
    .D(_00982_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[0] ));
 sky130_fd_sc_hd__dfxtp_1 _24450_ (.CLK(clknet_leaf_64_clk),
    .D(_00983_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24451_ (.CLK(clknet_leaf_63_clk),
    .D(_00984_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[2] ));
 sky130_fd_sc_hd__dfxtp_1 _24452_ (.CLK(clknet_leaf_64_clk),
    .D(_00985_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[3] ));
 sky130_fd_sc_hd__dfxtp_1 _24453_ (.CLK(clknet_leaf_62_clk),
    .D(_00986_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24454_ (.CLK(clknet_leaf_62_clk),
    .D(_00987_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[5] ));
 sky130_fd_sc_hd__dfxtp_2 _24455_ (.CLK(clknet_leaf_54_clk),
    .D(_00988_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24456_ (.CLK(clknet_4_15__leaf_clk),
    .D(_00989_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24457_ (.CLK(clknet_leaf_58_clk),
    .D(_00990_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[8] ));
 sky130_fd_sc_hd__dfxtp_1 _24458_ (.CLK(clknet_leaf_52_clk),
    .D(_00991_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[9] ));
 sky130_fd_sc_hd__dfxtp_1 _24459_ (.CLK(clknet_leaf_54_clk),
    .D(_00992_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[10] ));
 sky130_fd_sc_hd__dfxtp_1 _24460_ (.CLK(clknet_leaf_55_clk),
    .D(_00993_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[11] ));
 sky130_fd_sc_hd__dfxtp_1 _24461_ (.CLK(clknet_leaf_55_clk),
    .D(_00994_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[12] ));
 sky130_fd_sc_hd__dfxtp_1 _24462_ (.CLK(clknet_leaf_57_clk),
    .D(_00995_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[13] ));
 sky130_fd_sc_hd__dfxtp_1 _24463_ (.CLK(clknet_leaf_59_clk),
    .D(_00996_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[14] ));
 sky130_fd_sc_hd__dfxtp_1 _24464_ (.CLK(clknet_leaf_54_clk),
    .D(_00997_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[15] ));
 sky130_fd_sc_hd__dfxtp_1 _24465_ (.CLK(clknet_leaf_57_clk),
    .D(_00998_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[16] ));
 sky130_fd_sc_hd__dfxtp_1 _24466_ (.CLK(clknet_leaf_57_clk),
    .D(_00999_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[17] ));
 sky130_fd_sc_hd__dfxtp_1 _24467_ (.CLK(clknet_leaf_55_clk),
    .D(_01000_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[18] ));
 sky130_fd_sc_hd__dfxtp_1 _24468_ (.CLK(clknet_leaf_54_clk),
    .D(_01001_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[19] ));
 sky130_fd_sc_hd__dfxtp_1 _24469_ (.CLK(clknet_leaf_40_clk),
    .D(_01002_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[20] ));
 sky130_fd_sc_hd__dfxtp_1 _24470_ (.CLK(clknet_leaf_55_clk),
    .D(_01003_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[21] ));
 sky130_fd_sc_hd__dfxtp_1 _24471_ (.CLK(clknet_leaf_37_clk),
    .D(_01004_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[22] ));
 sky130_fd_sc_hd__dfxtp_1 _24472_ (.CLK(clknet_leaf_55_clk),
    .D(_01005_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[23] ));
 sky130_fd_sc_hd__dfxtp_1 _24473_ (.CLK(clknet_leaf_37_clk),
    .D(_01006_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[24] ));
 sky130_fd_sc_hd__dfxtp_1 _24474_ (.CLK(clknet_leaf_37_clk),
    .D(_01007_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[25] ));
 sky130_fd_sc_hd__dfxtp_1 _24475_ (.CLK(clknet_leaf_37_clk),
    .D(_01008_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[26] ));
 sky130_fd_sc_hd__dfxtp_1 _24476_ (.CLK(clknet_leaf_39_clk),
    .D(_01009_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[27] ));
 sky130_fd_sc_hd__dfxtp_1 _24477_ (.CLK(clknet_leaf_38_clk),
    .D(_01010_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[28] ));
 sky130_fd_sc_hd__dfxtp_1 _24478_ (.CLK(clknet_leaf_37_clk),
    .D(_01011_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[29] ));
 sky130_fd_sc_hd__dfxtp_1 _24479_ (.CLK(clknet_leaf_55_clk),
    .D(_01012_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[30] ));
 sky130_fd_sc_hd__dfxtp_1 _24480_ (.CLK(clknet_leaf_55_clk),
    .D(_01013_),
    .Q(\top_inst.axis_in_inst.inbuf_bus[31] ));
 sky130_fd_sc_hd__dfxtp_4 _24481_ (.CLK(clknet_leaf_46_clk),
    .D(_01014_),
    .Q(\top_inst.axis_in_inst.inbuf_valid ));
 sky130_fd_sc_hd__dfxtp_1 _24482_ (.CLK(clknet_leaf_115_clk),
    .D(_01015_),
    .Q(\top_inst.valid_pipe[0] ));
 sky130_fd_sc_hd__dfxtp_1 _24483_ (.CLK(clknet_leaf_115_clk),
    .D(_01016_),
    .Q(\top_inst.valid_pipe[1] ));
 sky130_fd_sc_hd__dfxtp_1 _24484_ (.CLK(clknet_leaf_115_clk),
    .D(_01017_),
    .Q(\top_inst.valid_pipe[2] ));
 sky130_fd_sc_hd__dfxtp_1 _24485_ (.CLK(clknet_leaf_115_clk),
    .D(_01018_),
    .Q(\top_inst.valid_pipe[3] ));
 sky130_fd_sc_hd__dfxtp_1 _24486_ (.CLK(clknet_leaf_84_clk),
    .D(net285),
    .Q(\top_inst.valid_pipe[4] ));
 sky130_fd_sc_hd__dfxtp_1 _24487_ (.CLK(clknet_leaf_84_clk),
    .D(_01020_),
    .Q(\top_inst.valid_pipe[5] ));
 sky130_fd_sc_hd__dfxtp_1 _24488_ (.CLK(clknet_leaf_15_clk),
    .D(_01021_),
    .Q(\top_inst.valid_pipe[6] ));
 sky130_fd_sc_hd__dfxtp_1 _24489_ (.CLK(clknet_leaf_45_clk),
    .D(net332),
    .Q(\top_inst.valid_pipe[7] ));
 sky130_fd_sc_hd__dfxtp_1 _24490_ (.CLK(clknet_leaf_45_clk),
    .D(_01023_),
    .Q(\top_inst.axis_out_inst.out_buff_enabled ));
 sky130_fd_sc_hd__dfxtp_4 _24491_ (.CLK(clknet_leaf_109_clk),
    .D(_01024_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_2 _24492_ (.CLK(clknet_leaf_109_clk),
    .D(_01025_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_4 _24493_ (.CLK(clknet_leaf_125_clk),
    .D(_01026_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_2 _24494_ (.CLK(clknet_leaf_108_clk),
    .D(_01027_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_4 _24495_ (.CLK(clknet_leaf_125_clk),
    .D(_01028_),
    .Q(net110));
 sky130_fd_sc_hd__dfxtp_2 _24496_ (.CLK(clknet_leaf_126_clk),
    .D(_01029_),
    .Q(net121));
 sky130_fd_sc_hd__dfxtp_2 _24497_ (.CLK(clknet_leaf_108_clk),
    .D(_01030_),
    .Q(net132));
 sky130_fd_sc_hd__dfxtp_4 _24498_ (.CLK(clknet_leaf_125_clk),
    .D(_01031_),
    .Q(net143));
 sky130_fd_sc_hd__dfxtp_4 _24499_ (.CLK(clknet_leaf_128_clk),
    .D(_01032_),
    .Q(net154));
 sky130_fd_sc_hd__dfxtp_2 _24500_ (.CLK(clknet_leaf_126_clk),
    .D(_01033_),
    .Q(net165));
 sky130_fd_sc_hd__dfxtp_4 _24501_ (.CLK(clknet_leaf_128_clk),
    .D(_01034_),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_4 _24502_ (.CLK(clknet_leaf_123_clk),
    .D(_01035_),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_4 _24503_ (.CLK(clknet_leaf_127_clk),
    .D(_01036_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_2 _24504_ (.CLK(clknet_leaf_128_clk),
    .D(_01037_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_4 _24505_ (.CLK(clknet_leaf_126_clk),
    .D(_01038_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_4 _24506_ (.CLK(clknet_leaf_128_clk),
    .D(_01039_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_2 _24507_ (.CLK(clknet_leaf_132_clk),
    .D(_01040_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_4 _24508_ (.CLK(clknet_leaf_127_clk),
    .D(_01041_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_4 _24509_ (.CLK(clknet_leaf_128_clk),
    .D(_01042_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_1 _24510_ (.CLK(clknet_leaf_128_clk),
    .D(_01043_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_4 _24511_ (.CLK(clknet_leaf_132_clk),
    .D(_01044_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_4 _24512_ (.CLK(clknet_leaf_135_clk),
    .D(_01045_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_1 _24513_ (.CLK(clknet_leaf_132_clk),
    .D(_01046_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_2 _24514_ (.CLK(clknet_leaf_132_clk),
    .D(_01047_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_4 _24515_ (.CLK(clknet_leaf_132_clk),
    .D(_01048_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_1 _24516_ (.CLK(clknet_leaf_133_clk),
    .D(_01049_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_4 _24517_ (.CLK(clknet_leaf_135_clk),
    .D(_01050_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_2 _24518_ (.CLK(clknet_leaf_135_clk),
    .D(_01051_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_4 _24519_ (.CLK(clknet_leaf_132_clk),
    .D(_01052_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_4 _24520_ (.CLK(clknet_leaf_132_clk),
    .D(_01053_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_4 _24521_ (.CLK(clknet_leaf_128_clk),
    .D(_01054_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_4 _24522_ (.CLK(clknet_leaf_131_clk),
    .D(_01055_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_4 _24523_ (.CLK(clknet_leaf_128_clk),
    .D(_01056_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_2 _24524_ (.CLK(clknet_leaf_131_clk),
    .D(_01057_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_4 _24525_ (.CLK(clknet_leaf_128_clk),
    .D(_01058_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_2 _24526_ (.CLK(clknet_leaf_128_clk),
    .D(_01059_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_4 _24527_ (.CLK(clknet_leaf_128_clk),
    .D(_01060_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_1 _24528_ (.CLK(clknet_leaf_130_clk),
    .D(_01061_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_2 _24529_ (.CLK(clknet_leaf_130_clk),
    .D(_01062_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_4 _24530_ (.CLK(clknet_leaf_129_clk),
    .D(_01063_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_4 _24531_ (.CLK(clknet_leaf_129_clk),
    .D(_01064_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_4 _24532_ (.CLK(clknet_leaf_103_clk),
    .D(_01065_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_2 _24533_ (.CLK(clknet_leaf_130_clk),
    .D(_01066_),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_2 _24534_ (.CLK(clknet_leaf_131_clk),
    .D(_01067_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_2 _24535_ (.CLK(clknet_leaf_131_clk),
    .D(_01068_),
    .Q(net104));
 sky130_fd_sc_hd__dfxtp_2 _24536_ (.CLK(clknet_leaf_102_clk),
    .D(_01069_),
    .Q(net105));
 sky130_fd_sc_hd__dfxtp_4 _24537_ (.CLK(clknet_leaf_129_clk),
    .D(_01070_),
    .Q(net106));
 sky130_fd_sc_hd__dfxtp_4 _24538_ (.CLK(clknet_leaf_101_clk),
    .D(_01071_),
    .Q(net107));
 sky130_fd_sc_hd__dfxtp_4 _24539_ (.CLK(clknet_leaf_130_clk),
    .D(_01072_),
    .Q(net108));
 sky130_fd_sc_hd__dfxtp_4 _24540_ (.CLK(clknet_leaf_102_clk),
    .D(_01073_),
    .Q(net109));
 sky130_fd_sc_hd__dfxtp_2 _24541_ (.CLK(clknet_leaf_102_clk),
    .D(_01074_),
    .Q(net111));
 sky130_fd_sc_hd__dfxtp_4 _24542_ (.CLK(clknet_leaf_100_clk),
    .D(_01075_),
    .Q(net112));
 sky130_fd_sc_hd__dfxtp_4 _24543_ (.CLK(clknet_leaf_130_clk),
    .D(_01076_),
    .Q(net113));
 sky130_fd_sc_hd__dfxtp_2 _24544_ (.CLK(clknet_leaf_100_clk),
    .D(_01077_),
    .Q(net114));
 sky130_fd_sc_hd__dfxtp_2 _24545_ (.CLK(clknet_leaf_100_clk),
    .D(_01078_),
    .Q(net115));
 sky130_fd_sc_hd__dfxtp_1 _24546_ (.CLK(clknet_leaf_103_clk),
    .D(_01079_),
    .Q(net116));
 sky130_fd_sc_hd__dfxtp_4 _24547_ (.CLK(clknet_leaf_100_clk),
    .D(_01080_),
    .Q(net117));
 sky130_fd_sc_hd__dfxtp_4 _24548_ (.CLK(clknet_leaf_100_clk),
    .D(_01081_),
    .Q(net118));
 sky130_fd_sc_hd__dfxtp_2 _24549_ (.CLK(clknet_leaf_131_clk),
    .D(_01082_),
    .Q(net119));
 sky130_fd_sc_hd__dfxtp_2 _24550_ (.CLK(clknet_leaf_100_clk),
    .D(_01083_),
    .Q(net120));
 sky130_fd_sc_hd__dfxtp_2 _24551_ (.CLK(clknet_leaf_103_clk),
    .D(_01084_),
    .Q(net122));
 sky130_fd_sc_hd__dfxtp_4 _24552_ (.CLK(clknet_leaf_133_clk),
    .D(_01085_),
    .Q(net123));
 sky130_fd_sc_hd__dfxtp_2 _24553_ (.CLK(clknet_leaf_103_clk),
    .D(_01086_),
    .Q(net124));
 sky130_fd_sc_hd__dfxtp_2 _24554_ (.CLK(clknet_leaf_133_clk),
    .D(_01087_),
    .Q(net125));
 sky130_fd_sc_hd__dfxtp_1 _24555_ (.CLK(clknet_leaf_133_clk),
    .D(_01088_),
    .Q(net126));
 sky130_fd_sc_hd__dfxtp_2 _24556_ (.CLK(clknet_leaf_136_clk),
    .D(_01089_),
    .Q(net127));
 sky130_fd_sc_hd__dfxtp_4 _24557_ (.CLK(clknet_leaf_135_clk),
    .D(_01090_),
    .Q(net128));
 sky130_fd_sc_hd__dfxtp_4 _24558_ (.CLK(clknet_leaf_135_clk),
    .D(_01091_),
    .Q(net129));
 sky130_fd_sc_hd__dfxtp_4 _24559_ (.CLK(clknet_leaf_133_clk),
    .D(_01092_),
    .Q(net130));
 sky130_fd_sc_hd__dfxtp_2 _24560_ (.CLK(clknet_leaf_134_clk),
    .D(_01093_),
    .Q(net131));
 sky130_fd_sc_hd__dfxtp_4 _24561_ (.CLK(clknet_leaf_137_clk),
    .D(_01094_),
    .Q(net133));
 sky130_fd_sc_hd__dfxtp_4 _24562_ (.CLK(clknet_leaf_137_clk),
    .D(_01095_),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_4 _24563_ (.CLK(clknet_leaf_137_clk),
    .D(_01096_),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_4 _24564_ (.CLK(clknet_leaf_134_clk),
    .D(_01097_),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_4 _24565_ (.CLK(clknet_leaf_137_clk),
    .D(_01098_),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_4 _24566_ (.CLK(clknet_leaf_137_clk),
    .D(_01099_),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_4 _24567_ (.CLK(clknet_leaf_138_clk),
    .D(_01100_),
    .Q(net139));
 sky130_fd_sc_hd__dfxtp_2 _24568_ (.CLK(clknet_leaf_134_clk),
    .D(_01101_),
    .Q(net140));
 sky130_fd_sc_hd__dfxtp_2 _24569_ (.CLK(clknet_leaf_141_clk),
    .D(_01102_),
    .Q(net141));
 sky130_fd_sc_hd__dfxtp_2 _24570_ (.CLK(clknet_leaf_134_clk),
    .D(_01103_),
    .Q(net142));
 sky130_fd_sc_hd__dfxtp_1 _24571_ (.CLK(clknet_leaf_143_clk),
    .D(_01104_),
    .Q(net144));
 sky130_fd_sc_hd__dfxtp_4 _24572_ (.CLK(clknet_leaf_140_clk),
    .D(_01105_),
    .Q(net145));
 sky130_fd_sc_hd__dfxtp_2 _24573_ (.CLK(clknet_leaf_139_clk),
    .D(_01106_),
    .Q(net146));
 sky130_fd_sc_hd__dfxtp_1 _24574_ (.CLK(clknet_leaf_142_clk),
    .D(_01107_),
    .Q(net147));
 sky130_fd_sc_hd__dfxtp_2 _24575_ (.CLK(clknet_leaf_142_clk),
    .D(_01108_),
    .Q(net148));
 sky130_fd_sc_hd__dfxtp_1 _24576_ (.CLK(clknet_leaf_142_clk),
    .D(_01109_),
    .Q(net149));
 sky130_fd_sc_hd__dfxtp_4 _24577_ (.CLK(clknet_leaf_140_clk),
    .D(_01110_),
    .Q(net150));
 sky130_fd_sc_hd__dfxtp_2 _24578_ (.CLK(clknet_leaf_142_clk),
    .D(_01111_),
    .Q(net151));
 sky130_fd_sc_hd__dfxtp_4 _24579_ (.CLK(clknet_leaf_140_clk),
    .D(_01112_),
    .Q(net152));
 sky130_fd_sc_hd__dfxtp_4 _24580_ (.CLK(clknet_leaf_142_clk),
    .D(_01113_),
    .Q(net153));
 sky130_fd_sc_hd__dfxtp_1 _24581_ (.CLK(clknet_leaf_139_clk),
    .D(_01114_),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_1 _24582_ (.CLK(clknet_leaf_142_clk),
    .D(_01115_),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_1 _24583_ (.CLK(clknet_leaf_142_clk),
    .D(_01116_),
    .Q(net157));
 sky130_fd_sc_hd__dfxtp_1 _24584_ (.CLK(clknet_leaf_141_clk),
    .D(_01117_),
    .Q(net158));
 sky130_fd_sc_hd__dfxtp_4 _24585_ (.CLK(clknet_leaf_20_clk),
    .D(_01118_),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_2 _24586_ (.CLK(clknet_leaf_141_clk),
    .D(_01119_),
    .Q(net160));
 sky130_fd_sc_hd__dfxtp_4 _24587_ (.CLK(clknet_leaf_20_clk),
    .D(_01120_),
    .Q(net161));
 sky130_fd_sc_hd__dfxtp_4 _24588_ (.CLK(clknet_leaf_32_clk),
    .D(_01121_),
    .Q(net162));
 sky130_fd_sc_hd__dfxtp_2 _24589_ (.CLK(clknet_leaf_32_clk),
    .D(_01122_),
    .Q(net163));
 sky130_fd_sc_hd__dfxtp_2 _24590_ (.CLK(clknet_leaf_32_clk),
    .D(_01123_),
    .Q(net164));
 sky130_fd_sc_hd__dfxtp_2 _24591_ (.CLK(clknet_leaf_22_clk),
    .D(_01124_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_2 _24592_ (.CLK(clknet_leaf_22_clk),
    .D(_01125_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_2 _24593_ (.CLK(clknet_leaf_24_clk),
    .D(_01126_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_2 _24594_ (.CLK(clknet_leaf_22_clk),
    .D(_01127_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_4 _24595_ (.CLK(clknet_leaf_23_clk),
    .D(_01128_),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_2 _24596_ (.CLK(clknet_leaf_22_clk),
    .D(_01129_),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_4 _24597_ (.CLK(clknet_leaf_22_clk),
    .D(_01130_),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_4 _24598_ (.CLK(clknet_leaf_22_clk),
    .D(_01131_),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_4 _24599_ (.CLK(clknet_leaf_23_clk),
    .D(_01132_),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_2 _24600_ (.CLK(clknet_leaf_24_clk),
    .D(_01133_),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_2 _24601_ (.CLK(clknet_leaf_24_clk),
    .D(_01134_),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_4 _24602_ (.CLK(clknet_leaf_23_clk),
    .D(_01135_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_2 _24603_ (.CLK(clknet_leaf_30_clk),
    .D(_01136_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _24604_ (.CLK(clknet_leaf_21_clk),
    .D(_01137_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_4 _24605_ (.CLK(clknet_leaf_21_clk),
    .D(_01138_),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_4 _24606_ (.CLK(clknet_leaf_25_clk),
    .D(_01139_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_4 _24607_ (.CLK(clknet_leaf_25_clk),
    .D(_01140_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_4 _24608_ (.CLK(clknet_leaf_22_clk),
    .D(_01141_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_4 _24609_ (.CLK(clknet_leaf_21_clk),
    .D(_01142_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_4 _24610_ (.CLK(clknet_leaf_21_clk),
    .D(_01143_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_2 _24611_ (.CLK(clknet_leaf_21_clk),
    .D(_01144_),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_2 _24612_ (.CLK(clknet_leaf_31_clk),
    .D(_01145_),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_4 _24613_ (.CLK(clknet_leaf_21_clk),
    .D(_01146_),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_4 _24614_ (.CLK(clknet_leaf_21_clk),
    .D(_01147_),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_4 _24615_ (.CLK(clknet_leaf_32_clk),
    .D(_01148_),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_2 _24616_ (.CLK(clknet_leaf_31_clk),
    .D(_01149_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_4 _24617_ (.CLK(clknet_leaf_32_clk),
    .D(_01150_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_4 _24618_ (.CLK(clknet_leaf_21_clk),
    .D(_01151_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_4 _24619_ (.CLK(clknet_leaf_16_clk),
    .D(_01152_),
    .Q(net166));
 sky130_fd_sc_hd__dfxtp_1 _24620_ (.CLK(clknet_leaf_32_clk),
    .D(_01153_),
    .Q(\top_inst.axis_out_inst.out_buff_data[96] ));
 sky130_fd_sc_hd__dfxtp_1 _24621_ (.CLK(clknet_leaf_21_clk),
    .D(net582),
    .Q(\top_inst.axis_out_inst.out_buff_data[97] ));
 sky130_fd_sc_hd__dfxtp_1 _24622_ (.CLK(clknet_leaf_22_clk),
    .D(net532),
    .Q(\top_inst.axis_out_inst.out_buff_data[98] ));
 sky130_fd_sc_hd__dfxtp_1 _24623_ (.CLK(clknet_leaf_23_clk),
    .D(_01156_),
    .Q(\top_inst.axis_out_inst.out_buff_data[99] ));
 sky130_fd_sc_hd__dfxtp_1 _24624_ (.CLK(clknet_leaf_25_clk),
    .D(net372),
    .Q(\top_inst.axis_out_inst.out_buff_data[100] ));
 sky130_fd_sc_hd__dfxtp_1 _24625_ (.CLK(clknet_leaf_25_clk),
    .D(net425),
    .Q(\top_inst.axis_out_inst.out_buff_data[101] ));
 sky130_fd_sc_hd__dfxtp_1 _24626_ (.CLK(clknet_leaf_24_clk),
    .D(net303),
    .Q(\top_inst.axis_out_inst.out_buff_data[102] ));
 sky130_fd_sc_hd__dfxtp_1 _24627_ (.CLK(clknet_leaf_23_clk),
    .D(net291),
    .Q(\top_inst.axis_out_inst.out_buff_data[103] ));
 sky130_fd_sc_hd__dfxtp_1 _24628_ (.CLK(clknet_leaf_24_clk),
    .D(_01161_),
    .Q(\top_inst.axis_out_inst.out_buff_data[104] ));
 sky130_fd_sc_hd__dfxtp_1 _24629_ (.CLK(clknet_leaf_22_clk),
    .D(_01162_),
    .Q(\top_inst.axis_out_inst.out_buff_data[105] ));
 sky130_fd_sc_hd__dfxtp_1 _24630_ (.CLK(clknet_leaf_25_clk),
    .D(_01163_),
    .Q(\top_inst.axis_out_inst.out_buff_data[106] ));
 sky130_fd_sc_hd__dfxtp_1 _24631_ (.CLK(clknet_leaf_25_clk),
    .D(_01164_),
    .Q(\top_inst.axis_out_inst.out_buff_data[107] ));
 sky130_fd_sc_hd__dfxtp_1 _24632_ (.CLK(clknet_leaf_23_clk),
    .D(net660),
    .Q(\top_inst.axis_out_inst.out_buff_data[108] ));
 sky130_fd_sc_hd__dfxtp_1 _24633_ (.CLK(clknet_leaf_24_clk),
    .D(net628),
    .Q(\top_inst.axis_out_inst.out_buff_data[109] ));
 sky130_fd_sc_hd__dfxtp_1 _24634_ (.CLK(clknet_leaf_26_clk),
    .D(_01167_),
    .Q(\top_inst.axis_out_inst.out_buff_data[110] ));
 sky130_fd_sc_hd__dfxtp_1 _24635_ (.CLK(clknet_leaf_24_clk),
    .D(_01168_),
    .Q(\top_inst.axis_out_inst.out_buff_data[111] ));
 sky130_fd_sc_hd__dfxtp_1 _24636_ (.CLK(clknet_leaf_25_clk),
    .D(net509),
    .Q(\top_inst.axis_out_inst.out_buff_data[112] ));
 sky130_fd_sc_hd__dfxtp_1 _24637_ (.CLK(clknet_leaf_26_clk),
    .D(_01170_),
    .Q(\top_inst.axis_out_inst.out_buff_data[113] ));
 sky130_fd_sc_hd__dfxtp_1 _24638_ (.CLK(clknet_leaf_21_clk),
    .D(_01171_),
    .Q(\top_inst.axis_out_inst.out_buff_data[114] ));
 sky130_fd_sc_hd__dfxtp_1 _24639_ (.CLK(clknet_leaf_25_clk),
    .D(net543),
    .Q(\top_inst.axis_out_inst.out_buff_data[115] ));
 sky130_fd_sc_hd__dfxtp_1 _24640_ (.CLK(clknet_leaf_25_clk),
    .D(net534),
    .Q(\top_inst.axis_out_inst.out_buff_data[116] ));
 sky130_fd_sc_hd__dfxtp_1 _24641_ (.CLK(clknet_leaf_22_clk),
    .D(net261),
    .Q(\top_inst.axis_out_inst.out_buff_data[117] ));
 sky130_fd_sc_hd__dfxtp_1 _24642_ (.CLK(clknet_leaf_30_clk),
    .D(_01175_),
    .Q(\top_inst.axis_out_inst.out_buff_data[118] ));
 sky130_fd_sc_hd__dfxtp_1 _24643_ (.CLK(clknet_leaf_21_clk),
    .D(net609),
    .Q(\top_inst.axis_out_inst.out_buff_data[119] ));
 sky130_fd_sc_hd__dfxtp_1 _24644_ (.CLK(clknet_leaf_21_clk),
    .D(net442),
    .Q(\top_inst.axis_out_inst.out_buff_data[120] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(input_tdata[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input2 (.A(input_tdata[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(input_tdata[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(input_tdata[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(input_tdata[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(input_tdata[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(input_tdata[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(input_tdata[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(input_tdata[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 input10 (.A(input_tdata[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(input_tdata[19]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(input_tdata[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(input_tdata[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(input_tdata[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(input_tdata[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_4 input16 (.A(input_tdata[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(input_tdata[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input18 (.A(input_tdata[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(input_tdata[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(input_tdata[27]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(input_tdata[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(input_tdata[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_8 input23 (.A(input_tdata[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_8 input24 (.A(input_tdata[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_4 input25 (.A(input_tdata[31]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(input_tdata[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_8 input27 (.A(input_tdata[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(input_tdata[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(input_tdata[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(input_tdata[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(input_tdata[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(input_tdata[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_4 input33 (.A(input_tvalid),
    .X(net33));
 sky130_fd_sc_hd__buf_12 input34 (.A(load_weight),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(output_tready),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(reset),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 output37 (.A(net37),
    .X(input_tready));
 sky130_fd_sc_hd__clkbuf_4 output38 (.A(net38),
    .X(output_tdata[0]));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net39),
    .X(output_tdata[100]));
 sky130_fd_sc_hd__clkbuf_4 output40 (.A(net40),
    .X(output_tdata[101]));
 sky130_fd_sc_hd__clkbuf_4 output41 (.A(net41),
    .X(output_tdata[102]));
 sky130_fd_sc_hd__clkbuf_4 output42 (.A(net42),
    .X(output_tdata[103]));
 sky130_fd_sc_hd__clkbuf_4 output43 (.A(net43),
    .X(output_tdata[104]));
 sky130_fd_sc_hd__clkbuf_4 output44 (.A(net44),
    .X(output_tdata[105]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(output_tdata[106]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(output_tdata[107]));
 sky130_fd_sc_hd__clkbuf_4 output47 (.A(net47),
    .X(output_tdata[108]));
 sky130_fd_sc_hd__clkbuf_4 output48 (.A(net48),
    .X(output_tdata[109]));
 sky130_fd_sc_hd__clkbuf_4 output49 (.A(net49),
    .X(output_tdata[10]));
 sky130_fd_sc_hd__clkbuf_4 output50 (.A(net50),
    .X(output_tdata[110]));
 sky130_fd_sc_hd__clkbuf_4 output51 (.A(net51),
    .X(output_tdata[111]));
 sky130_fd_sc_hd__clkbuf_4 output52 (.A(net52),
    .X(output_tdata[112]));
 sky130_fd_sc_hd__clkbuf_4 output53 (.A(net53),
    .X(output_tdata[113]));
 sky130_fd_sc_hd__clkbuf_4 output54 (.A(net54),
    .X(output_tdata[114]));
 sky130_fd_sc_hd__clkbuf_4 output55 (.A(net55),
    .X(output_tdata[115]));
 sky130_fd_sc_hd__clkbuf_4 output56 (.A(net56),
    .X(output_tdata[116]));
 sky130_fd_sc_hd__clkbuf_4 output57 (.A(net57),
    .X(output_tdata[117]));
 sky130_fd_sc_hd__clkbuf_4 output58 (.A(net58),
    .X(output_tdata[118]));
 sky130_fd_sc_hd__clkbuf_4 output59 (.A(net59),
    .X(output_tdata[119]));
 sky130_fd_sc_hd__clkbuf_4 output60 (.A(net60),
    .X(output_tdata[11]));
 sky130_fd_sc_hd__clkbuf_4 output61 (.A(net61),
    .X(output_tdata[120]));
 sky130_fd_sc_hd__clkbuf_4 output62 (.A(net62),
    .X(output_tdata[121]));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net63),
    .X(output_tdata[122]));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net64),
    .X(output_tdata[123]));
 sky130_fd_sc_hd__clkbuf_4 output65 (.A(net65),
    .X(output_tdata[124]));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net66),
    .X(output_tdata[125]));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net67),
    .X(output_tdata[126]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(output_tdata[127]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(output_tdata[12]));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(output_tdata[13]));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net71),
    .X(output_tdata[14]));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .X(output_tdata[15]));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net73),
    .X(output_tdata[16]));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net74),
    .X(output_tdata[17]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(output_tdata[18]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(output_tdata[19]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(output_tdata[1]));
 sky130_fd_sc_hd__clkbuf_4 output78 (.A(net78),
    .X(output_tdata[20]));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net79),
    .X(output_tdata[21]));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net80),
    .X(output_tdata[22]));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net81),
    .X(output_tdata[23]));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net82),
    .X(output_tdata[24]));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net83),
    .X(output_tdata[25]));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net84),
    .X(output_tdata[26]));
 sky130_fd_sc_hd__clkbuf_4 output85 (.A(net85),
    .X(output_tdata[27]));
 sky130_fd_sc_hd__clkbuf_4 output86 (.A(net86),
    .X(output_tdata[28]));
 sky130_fd_sc_hd__clkbuf_4 output87 (.A(net87),
    .X(output_tdata[29]));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net88),
    .X(output_tdata[2]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(output_tdata[30]));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net90),
    .X(output_tdata[31]));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net91),
    .X(output_tdata[32]));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net92),
    .X(output_tdata[33]));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net93),
    .X(output_tdata[34]));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net94),
    .X(output_tdata[35]));
 sky130_fd_sc_hd__clkbuf_4 output95 (.A(net95),
    .X(output_tdata[36]));
 sky130_fd_sc_hd__clkbuf_4 output96 (.A(net96),
    .X(output_tdata[37]));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net97),
    .X(output_tdata[38]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(output_tdata[39]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(output_tdata[3]));
 sky130_fd_sc_hd__clkbuf_4 output100 (.A(net100),
    .X(output_tdata[40]));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net101),
    .X(output_tdata[41]));
 sky130_fd_sc_hd__clkbuf_4 output102 (.A(net102),
    .X(output_tdata[42]));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net103),
    .X(output_tdata[43]));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net104),
    .X(output_tdata[44]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(output_tdata[45]));
 sky130_fd_sc_hd__clkbuf_4 output106 (.A(net106),
    .X(output_tdata[46]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(output_tdata[47]));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net108),
    .X(output_tdata[48]));
 sky130_fd_sc_hd__clkbuf_4 output109 (.A(net109),
    .X(output_tdata[49]));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net110),
    .X(output_tdata[4]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(output_tdata[50]));
 sky130_fd_sc_hd__clkbuf_4 output112 (.A(net112),
    .X(output_tdata[51]));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net113),
    .X(output_tdata[52]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(output_tdata[53]));
 sky130_fd_sc_hd__clkbuf_4 output115 (.A(net115),
    .X(output_tdata[54]));
 sky130_fd_sc_hd__clkbuf_4 output116 (.A(net116),
    .X(output_tdata[55]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(output_tdata[56]));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net118),
    .X(output_tdata[57]));
 sky130_fd_sc_hd__clkbuf_4 output119 (.A(net119),
    .X(output_tdata[58]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(output_tdata[59]));
 sky130_fd_sc_hd__clkbuf_4 output121 (.A(net121),
    .X(output_tdata[5]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(output_tdata[60]));
 sky130_fd_sc_hd__clkbuf_4 output123 (.A(net123),
    .X(output_tdata[61]));
 sky130_fd_sc_hd__clkbuf_4 output124 (.A(net124),
    .X(output_tdata[62]));
 sky130_fd_sc_hd__clkbuf_4 output125 (.A(net125),
    .X(output_tdata[63]));
 sky130_fd_sc_hd__clkbuf_4 output126 (.A(net126),
    .X(output_tdata[64]));
 sky130_fd_sc_hd__clkbuf_4 output127 (.A(net127),
    .X(output_tdata[65]));
 sky130_fd_sc_hd__clkbuf_4 output128 (.A(net128),
    .X(output_tdata[66]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(output_tdata[67]));
 sky130_fd_sc_hd__clkbuf_4 output130 (.A(net130),
    .X(output_tdata[68]));
 sky130_fd_sc_hd__clkbuf_4 output131 (.A(net131),
    .X(output_tdata[69]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(output_tdata[6]));
 sky130_fd_sc_hd__clkbuf_4 output133 (.A(net133),
    .X(output_tdata[70]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(output_tdata[71]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(output_tdata[72]));
 sky130_fd_sc_hd__clkbuf_4 output136 (.A(net136),
    .X(output_tdata[73]));
 sky130_fd_sc_hd__clkbuf_4 output137 (.A(net137),
    .X(output_tdata[74]));
 sky130_fd_sc_hd__clkbuf_4 output138 (.A(net138),
    .X(output_tdata[75]));
 sky130_fd_sc_hd__clkbuf_4 output139 (.A(net139),
    .X(output_tdata[76]));
 sky130_fd_sc_hd__clkbuf_4 output140 (.A(net140),
    .X(output_tdata[77]));
 sky130_fd_sc_hd__clkbuf_4 output141 (.A(net141),
    .X(output_tdata[78]));
 sky130_fd_sc_hd__clkbuf_4 output142 (.A(net142),
    .X(output_tdata[79]));
 sky130_fd_sc_hd__clkbuf_4 output143 (.A(net143),
    .X(output_tdata[7]));
 sky130_fd_sc_hd__clkbuf_4 output144 (.A(net144),
    .X(output_tdata[80]));
 sky130_fd_sc_hd__clkbuf_4 output145 (.A(net145),
    .X(output_tdata[81]));
 sky130_fd_sc_hd__clkbuf_4 output146 (.A(net146),
    .X(output_tdata[82]));
 sky130_fd_sc_hd__clkbuf_4 output147 (.A(net147),
    .X(output_tdata[83]));
 sky130_fd_sc_hd__clkbuf_4 output148 (.A(net148),
    .X(output_tdata[84]));
 sky130_fd_sc_hd__clkbuf_4 output149 (.A(net149),
    .X(output_tdata[85]));
 sky130_fd_sc_hd__clkbuf_4 output150 (.A(net150),
    .X(output_tdata[86]));
 sky130_fd_sc_hd__clkbuf_4 output151 (.A(net151),
    .X(output_tdata[87]));
 sky130_fd_sc_hd__clkbuf_4 output152 (.A(net152),
    .X(output_tdata[88]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(output_tdata[89]));
 sky130_fd_sc_hd__clkbuf_4 output154 (.A(net154),
    .X(output_tdata[8]));
 sky130_fd_sc_hd__clkbuf_4 output155 (.A(net155),
    .X(output_tdata[90]));
 sky130_fd_sc_hd__clkbuf_4 output156 (.A(net156),
    .X(output_tdata[91]));
 sky130_fd_sc_hd__clkbuf_4 output157 (.A(net157),
    .X(output_tdata[92]));
 sky130_fd_sc_hd__clkbuf_4 output158 (.A(net158),
    .X(output_tdata[93]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(output_tdata[94]));
 sky130_fd_sc_hd__clkbuf_4 output160 (.A(net160),
    .X(output_tdata[95]));
 sky130_fd_sc_hd__clkbuf_4 output161 (.A(net161),
    .X(output_tdata[96]));
 sky130_fd_sc_hd__clkbuf_4 output162 (.A(net162),
    .X(output_tdata[97]));
 sky130_fd_sc_hd__clkbuf_4 output163 (.A(net163),
    .X(output_tdata[98]));
 sky130_fd_sc_hd__clkbuf_4 output164 (.A(net164),
    .X(output_tdata[99]));
 sky130_fd_sc_hd__clkbuf_4 output165 (.A(net165),
    .X(output_tdata[9]));
 sky130_fd_sc_hd__clkbuf_4 output166 (.A(net166),
    .X(output_tvalid));
 sky130_fd_sc_hd__buf_4 wire167 (.A(_11129_),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 max_cap168 (.A(_01790_),
    .X(net168));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire169 (.A(_05879_),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 max_cap170 (.A(_09313_),
    .X(net170));
 sky130_fd_sc_hd__buf_1 max_cap171 (.A(_07180_),
    .X(net171));
 sky130_fd_sc_hd__buf_1 max_cap172 (.A(_11720_),
    .X(net172));
 sky130_fd_sc_hd__buf_1 max_cap173 (.A(_07101_),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 max_cap174 (.A(_02360_),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 max_cap175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 max_cap176 (.A(_02320_),
    .X(net176));
 sky130_fd_sc_hd__buf_1 max_cap177 (.A(_02279_),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 max_cap178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 max_cap179 (.A(_02233_),
    .X(net179));
 sky130_fd_sc_hd__buf_1 max_cap180 (.A(_06934_),
    .X(net180));
 sky130_fd_sc_hd__buf_1 max_cap181 (.A(_06494_),
    .X(net181));
 sky130_fd_sc_hd__buf_1 max_cap182 (.A(_06052_),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_8__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_10__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_11__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_12__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_15__leaf_clk));
 sky130_fd_sc_hd__buf_1 rebuffer1 (.A(_09446_),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 rebuffer2 (.A(_05265_),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 rebuffer3 (.A(_05265_),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 rebuffer4 (.A(_05265_),
    .X(net186));
 sky130_fd_sc_hd__buf_1 rebuffer5 (.A(net186),
    .X(net187));
 sky130_fd_sc_hd__buf_8 split6 (.A(_05265_),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 rebuffer7 (.A(_11681_),
    .X(net189));
 sky130_fd_sc_hd__buf_6 rebuffer8 (.A(net189),
    .X(net190));
 sky130_fd_sc_hd__buf_1 rebuffer9 (.A(net190),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 rebuffer10 (.A(net190),
    .X(net192));
 sky130_fd_sc_hd__buf_6 rebuffer11 (.A(_11699_),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 rebuffer12 (.A(net193),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 rebuffer13 (.A(net194),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 rebuffer14 (.A(_01458_),
    .X(net196));
 sky130_fd_sc_hd__buf_1 rebuffer15 (.A(_01266_),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 rebuffer16 (.A(net197),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 rebuffer17 (.A(_09721_),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 rebuffer18 (.A(_09464_),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 rebuffer19 (.A(_09519_),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 rebuffer20 (.A(_09214_),
    .X(net202));
 sky130_fd_sc_hd__buf_6 rebuffer21 (.A(_09214_),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 rebuffer22 (.A(_09518_),
    .X(net204));
 sky130_fd_sc_hd__buf_1 rebuffer23 (.A(_07059_),
    .X(net205));
 sky130_fd_sc_hd__buf_4 rebuffer24 (.A(_07059_),
    .X(net206));
 sky130_fd_sc_hd__buf_1 rebuffer25 (.A(net206),
    .X(net207));
 sky130_fd_sc_hd__buf_6 rebuffer26 (.A(net206),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 rebuffer27 (.A(_07167_),
    .X(net209));
 sky130_fd_sc_hd__buf_1 rebuffer28 (.A(_01384_),
    .X(net210));
 sky130_fd_sc_hd__buf_4 rebuffer29 (.A(_05266_),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 rebuffer30 (.A(net211),
    .X(net212));
 sky130_fd_sc_hd__buf_1 rebuffer31 (.A(net211),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 rebuffer32 (.A(_09522_),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 rebuffer33 (.A(_09205_),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 rebuffer34 (.A(_09205_),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_1 rebuffer35 (.A(net216),
    .X(net217));
 sky130_fd_sc_hd__buf_1 rebuffer36 (.A(_01234_),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 split37 (.A(_09218_),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_1 rebuffer38 (.A(_09514_),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_1 rebuffer39 (.A(_09555_),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_1 rebuffer40 (.A(net221),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_1 rebuffer41 (.A(_09196_),
    .X(net223));
 sky130_fd_sc_hd__buf_1 rebuffer42 (.A(_09196_),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 rebuffer43 (.A(net224),
    .X(net225));
 sky130_fd_sc_hd__buf_1 rebuffer44 (.A(_09517_),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 rebuffer45 (.A(_09205_),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 rebuffer46 (.A(_02827_),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_2 split47 (.A(_07593_),
    .X(net229));
 sky130_fd_sc_hd__buf_1 rebuffer48 (.A(_07196_),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_1 rebuffer49 (.A(_01262_),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_1 rebuffer50 (.A(_01266_),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 rebuffer51 (.A(net239),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 rebuffer52 (.A(net239),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 rebuffer53 (.A(_11699_),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 rebuffer54 (.A(_01282_),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_1 rebuffer55 (.A(_01285_),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 rebuffer56 (.A(_01462_),
    .X(net238));
 sky130_fd_sc_hd__buf_6 rebuffer57 (.A(_11691_),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 rebuffer58 (.A(net239),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 rebuffer59 (.A(_01330_),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_1 rebuffer60 (.A(_11676_),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_2 rebuffer61 (.A(net242),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 rebuffer62 (.A(net243),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_1 rebuffer63 (.A(net243),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_1 rebuffer64 (.A(_11686_),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 rebuffer65 (.A(net246),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_1 rebuffer66 (.A(net247),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 rebuffer67 (.A(_01401_),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 rebuffer68 (.A(_01501_),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 rebuffer69 (.A(net250),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][19] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_00154_),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][27] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_00162_),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\top_inst.axis_in_inst.inbuf_bus[7] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_00981_),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\top_inst.deskew_buff_inst.col_input[117] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_01174_),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][20] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_00155_),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][23] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_00158_),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][28] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_00163_),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\top_inst.deskew_buff_inst.col_input[50] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_00121_),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\top_inst.deskew_buff_inst.col_input[48] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_00119_),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][13] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_00148_),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][26] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_00161_),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][25] ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_00288_),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\top_inst.deskew_buff_inst.col_input[47] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_00118_),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\top_inst.deskew_buff_inst.col_input[49] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_00120_),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\top_inst.deskew_buff_inst.col_input[66] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_00041_),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\top_inst.valid_pipe[3] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_01019_),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][24] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_00287_),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][26] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_00289_),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\top_inst.deskew_buff_inst.col_input[103] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_01160_),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][20] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_00283_),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][6] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_00924_),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][3] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_00929_),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][21] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_00284_),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][31] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_00294_),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\top_inst.deskew_buff_inst.col_input[102] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_01159_),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][29] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_00292_),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][27] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_00258_),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][28] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_00195_),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\top_inst.axis_out_inst.out_buff_data[8] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\top_inst.deskew_buff_inst.col_input[16] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_00215_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\top_inst.deskew_buff_inst.col_input[67] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_00042_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\top_inst.deskew_buff_inst.col_input[46] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_00117_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\top_inst.axis_out_inst.out_buff_data[13] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\top_inst.deskew_buff_inst.col_input[99] ),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][17] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_00280_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][23] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_00286_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][15] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_00182_),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\top_inst.deskew_buff_inst.col_input[65] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_00040_),
    .X(net326));
 sky130_fd_sc_hd__buf_1 hold145 (.A(\top_inst.deskew_buff_inst.col_input[61] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_00132_),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][19] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_00282_),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\top_inst.valid_pipe[6] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_01022_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][22] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_00285_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][30] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_00293_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][7] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_00014_),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][30] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_00197_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][18] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_00185_),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\top_inst.deskew_buff_inst.col_input[3] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_00202_),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][18] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][16] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_00183_),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][4] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_00011_),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][19] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(_00186_),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][22] ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_00189_),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\top_inst.valid_pipe[5] ),
    .X(net354));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold173 (.A(\top_inst.deskew_buff_inst.col_input[4] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_00203_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][10] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_00177_),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\top_inst.axis_out_inst.out_buff_data[14] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][6] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_00013_),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][5] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_00012_),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\top_inst.axis_out_inst.out_buff_data[66] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][23] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_00190_),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][9] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_00016_),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][27] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_00290_),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\top_inst.deskew_buff_inst.col_input[100] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_01157_),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][9] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_00176_),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][29] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_00196_),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\top_inst.axis_out_inst.out_buff_data[67] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\top_inst.axis_out_inst.out_buff_data[36] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\top_inst.axis_out_inst.out_buff_data[24] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][6] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_00940_),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\top_inst.axis_out_inst.out_buff_data[20] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][31] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_00198_),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][24] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_00159_),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][2] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_00920_),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][5] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_00939_),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\top_inst.axis_out_inst.out_buff_data[85] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\top_inst.axis_out_inst.out_buff_data[113] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\top_inst.axis_out_inst.out_buff_data[84] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][6] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_00908_),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][0] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_00934_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][4] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_00171_),
    .X(net399));
 sky130_fd_sc_hd__buf_1 hold218 (.A(\top_inst.deskew_buff_inst.col_input[30] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_00229_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][6] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_00173_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][7] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_00957_),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][3] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_00905_),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\top_inst.deskew_buff_inst.col_input[2] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_00201_),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\top_inst.axis_out_inst.out_buff_data[123] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\top_inst.deskew_buff_inst.col_input[80] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_00055_),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][3] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_00937_),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\top_inst.axis_out_inst.out_buff_data[89] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][4] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_00938_),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][7] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_00174_),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\top_inst.deskew_buff_inst.col_input[11] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_00210_),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\top_inst.axis_out_inst.out_buff_data[4] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\top_inst.axis_out_inst.out_buff_data[110] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\top_inst.deskew_buff_inst.col_input[101] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(_01158_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\top_inst.deskew_buff_inst.col_input[10] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_00209_),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][31] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_00038_),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\top_inst.deskew_buff_inst.col_input[90] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_00065_),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][1] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_00168_),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\top_inst.axis_out_inst.out_buff_data[92] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\top_inst.deskew_buff_inst.col_input[18] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_00217_),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\top_inst.deskew_buff_inst.col_input[15] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(_00214_),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][12] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\top_inst.axis_out_inst.out_buff_data[10] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\top_inst.deskew_buff_inst.col_input[120] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_01177_),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\top_inst.axis_out_inst.out_buff_data[106] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\top_inst.axis_out_inst.out_buff_data[107] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][8] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_00143_),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][1] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_00136_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][12] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_00275_),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\top_inst.axis_out_inst.out_buff_data[122] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][5] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(_00268_),
    .X(net453));
 sky130_fd_sc_hd__buf_1 hold272 (.A(\top_inst.deskew_buff_inst.col_input[64] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_00039_),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][3] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(_00266_),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][6] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(_00141_),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\top_inst.axis_out_inst.out_buff_data[111] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\top_inst.axis_out_inst.out_buff_data[104] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\top_inst.axis_out_inst.out_buff_data[81] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\top_inst.axis_out_inst.out_buff_data[3] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\top_inst.deskew_buff_inst.col_input[9] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(_00208_),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][1] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\top_inst.axis_out_inst.out_buff_enabled ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\top_inst.axis_out_inst.out_buff_data[77] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][21] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_00156_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\top_inst.deskew_buff_inst.col_input[126] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_00005_),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\top_inst.axis_out_inst.out_buff_data[101] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][22] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_00029_),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\top_inst.axis_out_inst.out_buff_data[70] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\top_inst.deskew_buff_inst.col_input[58] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][3] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(_00074_),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][16] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][2] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_00073_),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\top_inst.deskew_buff_inst.col_input[14] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_00213_),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\top_inst.axis_out_inst.out_buff_data[17] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][18] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(_00153_),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][10] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\top_inst.axis_out_inst.out_buff_data[71] ),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_2 hold308 (.A(\top_inst.deskew_buff_inst.col_input[31] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(_00230_),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\top_inst.axis_out_inst.out_buff_data[30] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\top_inst.axis_out_inst.out_buff_data[32] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][3] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][0] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_00263_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\top_inst.deskew_buff_inst.col_input[36] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(_00107_),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\top_inst.deskew_buff_inst.col_input[127] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(_00006_),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][17] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_00152_),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\top_inst.deskew_buff_inst.col_input[82] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_00057_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][15] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][29] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(_00164_),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\top_inst.deskew_buff_inst.col_input[112] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(_01169_),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][22] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(_00157_),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\top_inst.axis_out_inst.out_buff_data[100] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\top_inst.axis_out_inst.out_buff_data[44] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][3] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][14] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(_00277_),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\top_inst.axis_out_inst.out_buff_data[118] ),
    .X(net517));
 sky130_fd_sc_hd__buf_1 hold336 (.A(\top_inst.deskew_buff_inst.col_input[63] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(_00134_),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][9] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(_00080_),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][18] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(_00025_),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\top_inst.deskew_buff_inst.col_input[88] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(_00063_),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][25] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(_00192_),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][7] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(_00238_),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\top_inst.axis_out_inst.out_buff_data[127] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\top_inst.deskew_buff_inst.col_input[98] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_01155_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\top_inst.deskew_buff_inst.col_input[116] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_01173_),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][11] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_00274_),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\top_inst.axis_out_inst.out_buff_data[82] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][14] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(_00149_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][21] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\top_inst.axis_out_inst.out_buff_data[6] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\top_inst.deskew_buff_inst.col_input[115] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(_01172_),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\top_inst.deskew_buff_inst.col_input[79] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(_00054_),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][7] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(_00142_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\top_inst.axis_out_inst.out_buff_data[25] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][13] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(_00084_),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][28] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_00099_),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\top_inst.axis_out_inst.out_buff_data[48] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][6] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(_00237_),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][2] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\top_inst.axis_out_inst.out_buff_data[95] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][4] ),
    .X(net558));
 sky130_fd_sc_hd__buf_1 hold377 (.A(\top_inst.deskew_buff_inst.col_input[62] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_00133_),
    .X(net560));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold379 (.A(\top_inst.deskew_buff_inst.col_input[93] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_00068_),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][11] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\top_inst.deskew_buff_inst.col_input[124] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(_00003_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][13] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][13] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][8] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(_00271_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][14] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(_00021_),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][9] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][16] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_00151_),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\top_inst.axis_out_inst.out_buff_data[98] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][17] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][9] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][1] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(_00903_),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\top_inst.valid_pipe[0] ),
    .X(net580));
 sky130_fd_sc_hd__buf_1 hold399 (.A(\top_inst.deskew_buff_inst.col_input[97] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_01154_),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\top_inst.axis_in_inst.inbuf_bus[14] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_00972_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\top_inst.deskew_buff_inst.col_input[7] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][17] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][15] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(_00150_),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][0] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\top_inst.axis_in_inst.inbuf_bus[20] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(_00946_),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][11] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(_00178_),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][3] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\top_inst.axis_out_inst.out_buff_data[40] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\top_inst.deskew_buff_inst.col_input[13] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(_00212_),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][29] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\top_inst.axis_out_inst.out_buff_data[91] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][4] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(_00235_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][1] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(_00959_),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\top_inst.deskew_buff_inst.col_input[68] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\top_inst.valid_pipe[2] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\top_inst.axis_in_inst.inbuf_bus[8] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(_00966_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\top_inst.deskew_buff_inst.col_input[119] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(_01176_),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\top_inst.axis_out_inst.out_buff_data[43] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\top_inst.deskew_buff_inst.col_input[78] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][5] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\top_inst.axis_out_inst.out_buff_data[42] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][15] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(_00022_),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\top_inst.axis_in_inst.inbuf_bus[5] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(_00979_),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\top_inst.axis_out_inst.out_buff_data[12] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\top_inst.axis_out_inst.out_buff_data[96] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\top_inst.valid_pipe[7] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][6] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\top_inst.axis_out_inst.out_buff_data[65] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\top_inst.axis_out_inst.out_buff_data[126] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\top_inst.valid_pipe[1] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][0] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_00007_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\top_inst.deskew_buff_inst.col_input[109] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(_01166_),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\top_inst.axis_out_inst.out_buff_data[87] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\top_inst.deskew_buff_inst.col_input[122] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\top_inst.deskew_buff_inst.col_input[42] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\top_inst.axis_out_inst.out_buff_data[11] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][7] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(_00965_),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\top_inst.axis_out_inst.out_buff_data[117] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\top_inst.deskew_buff_inst.col_input[86] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][6] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(_00964_),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[24] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][16] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(_00023_),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][1] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][1] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(_00951_),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\top_inst.axis_out_inst.out_buff_data[73] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[31] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\top_inst.deskew_buff_inst.col_input[55] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\top_inst.deskew_buff_inst.col_input[85] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(_00060_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][22] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\top_inst.axis_out_inst.out_buff_data[47] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][25] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\top_inst.valid_pipe[4] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\top_inst.deskew_buff_inst.col_input[111] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][2] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(_00904_),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\top_inst.axis_out_inst.out_buff_data[88] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\top_inst.axis_out_inst.out_buff_data[86] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\top_inst.deskew_buff_inst.col_input[108] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(_01165_),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\top_inst.axis_out_inst.out_buff_data[9] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][2] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(_00952_),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][30] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\top_inst.axis_out_inst.out_buff_data[39] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\top_inst.deskew_buff_inst.col_input[125] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(_00004_),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\top_inst.deskew_buff_inst.col_input[92] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(_00067_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\top_inst.deskew_buff_inst.col_input[87] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(_00062_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\top_inst.deskew_buff_inst.col_input[54] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\top_inst.axis_out_inst.out_buff_data[33] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][5] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(_00907_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\top_inst.axis_out_inst.out_buff_data[37] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\top_inst.axis_out_inst.out_buff_data[2] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][20] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\top_inst.axis_out_inst.out_buff_data[102] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][28] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][4] ),
    .X(net681));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold500 (.A(\top_inst.deskew_buff_inst.col_input[91] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(_00066_),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][29] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(_00036_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\top_inst.axis_out_inst.out_buff_data[5] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\top_inst.axis_out_inst.out_buff_data[79] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][27] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][30] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\top_inst.axis_out_inst.out_buff_data[69] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][28] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][14] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\top_inst.axis_out_inst.out_buff_data[51] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\top_inst.axis_out_inst.out_buff_data[90] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][29] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\top_inst.deskew_buff_inst.col_input[56] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\top_inst.axis_out_inst.out_buff_data[105] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][24] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\top_inst.axis_out_inst.out_buff_data[49] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][23] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(_00094_),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][3] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(_00961_),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][3] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\top_inst.axis_out_inst.out_buff_data[76] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[31] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][3] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][7] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(_00925_),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\top_inst.axis_out_inst.out_buff_data[112] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\top_inst.deskew_buff_inst.col_input[107] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][7] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(_00941_),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\top_inst.axis_out_inst.out_buff_data[109] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][0] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_00918_),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][0] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][4] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(_00962_),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][27] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(_00098_),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][31] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\top_inst.axis_out_inst.out_buff_data[26] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\top_inst.deskew_buff_inst.col_input[123] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\top_inst.axis_out_inst.out_buff_data[114] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][23] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\top_inst.axis_out_inst.out_buff_data[75] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][1] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\top_inst.axis_out_inst.out_buff_data[120] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(\top_inst.axis_out_inst.out_buff_data[62] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\top_inst.axis_out_inst.out_buff_data[46] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[0][0] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][15] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][0] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(_00958_),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\top_inst.axis_out_inst.out_buff_data[29] ),
    .X(net736));
 sky130_fd_sc_hd__buf_1 hold555 (.A(\top_inst.deskew_buff_inst.col_input[32] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_00103_),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\top_inst.axis_out_inst.out_buff_data[119] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\top_inst.deskew_buff_inst.col_input[114] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][5] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\top_inst.axis_out_inst.out_buff_data[83] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\top_inst.axis_out_inst.out_buff_data[74] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][1] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\top_inst.deskew_buff_inst.col_input[39] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][5] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][26] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[31] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\top_inst.axis_out_inst.out_buff_data[28] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][3] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\top_inst.axis_out_inst.out_buff_data[125] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\top_inst.axis_out_inst.out_buff_data[60] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\top_inst.deskew_buff_inst.col_input[75] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_00050_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\top_inst.axis_out_inst.out_buff_data[7] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\top_inst.deskew_buff_inst.col_input[28] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\top_inst.axis_out_inst.out_buff_data[72] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(\top_inst.deskew_buff_inst.col_input[35] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][20] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\top_inst.deskew_buff_inst.col_input[33] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][2] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][1] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\top_inst.axis_out_inst.out_buff_data[45] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][7] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(_00933_),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][2] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(_00936_),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\top_inst.axis_out_inst.out_buff_data[27] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\top_inst.skew_buff_inst.row[2].has_delay.shift_reg[1][1] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_00935_),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][6] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][2] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(_00960_),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\top_inst.axis_out_inst.out_buff_data[18] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][8] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\top_inst.axis_out_inst.out_buff_data[64] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\top_inst.deskew_buff_inst.col_input[121] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_00000_),
    .X(net778));
 sky130_fd_sc_hd__buf_1 hold597 (.A(\top_inst.deskew_buff_inst.col_input[34] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][4] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\top_inst.axis_out_inst.out_buff_data[97] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\top_inst.deskew_buff_inst.col_input[53] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][19] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][4] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(_00930_),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(\top_inst.deskew_buff_inst.col_input[24] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\top_inst.axis_out_inst.out_buff_data[1] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\top_inst.axis_out_inst.out_buff_data[116] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\top_inst.axis_out_inst.out_buff_data[34] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\top_inst.deskew_buff_inst.col_input[29] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][25] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(_00096_),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][25] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][26] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\top_inst.deskew_buff_inst.col_input[43] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(\top_inst.axis_out_inst.out_buff_data[50] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][5] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(_00140_),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\top_inst.axis_out_inst.out_buff_data[21] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][19] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\top_inst.axis_out_inst.out_buff_data[124] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(\top_inst.axis_out_inst.out_buff_data[54] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][8] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\top_inst.axis_out_inst.out_buff_data[78] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][21] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(_00092_),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][10] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\top_inst.deskew_buff_inst.col_input[72] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][4] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\top_inst.axis_out_inst.out_buff_data[115] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][18] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\top_inst.deskew_buff_inst.col_input[5] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(_00204_),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][24] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(_00095_),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\top_inst.deskew_buff_inst.col_input[44] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\top_inst.deskew_buff_inst.col_input[104] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\top_inst.deskew_buff_inst.col_input[77] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(_00052_),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][30] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\top_inst.axis_out_inst.out_buff_data[57] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\top_inst.axis_out_inst.out_buff_data[41] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][30] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][13] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\top_inst.deskew_buff_inst.col_input[22] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\top_inst.deskew_buff_inst.col_input[12] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(_00211_),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[0][5] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][11] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\top_inst.axis_out_inst.out_buff_data[19] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\top_inst.axis_out_inst.out_buff_data[93] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\top_inst.axis_out_inst.out_buff_data[16] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\top_inst.axis_out_inst.out_buff_data[108] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\top_inst.deskew_buff_inst.col_input[110] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][2] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][21] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\top_inst.deskew_buff_inst.col_input[45] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\top_inst.axis_out_inst.out_buff_data[56] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\top_inst.deskew_buff_inst.col_input[76] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(_00051_),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][10] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\top_inst.axis_out_inst.out_buff_data[121] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\top_inst.axis_out_inst.out_buff_data[23] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(\top_inst.axis_out_inst.out_buff_data[35] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\top_inst.axis_out_inst.out_buff_data[38] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(\top_inst.deskew_buff_inst.col_input[8] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(_00207_),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][2] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][22] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][7] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(_00909_),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[1][0] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(_00926_),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][31] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][12] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][13] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][12] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][2] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[27] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\top_inst.deskew_buff_inst.col_input[70] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\top_inst.deskew_buff_inst.col_input[52] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\top_inst.deskew_buff_inst.col_input[38] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][19] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][18] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][23] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][10] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[1] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\top_inst.deskew_buff_inst.col_input[94] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\top_inst.deskew_buff_inst.col_input[60] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\top_inst.axis_out_inst.out_buff_data[22] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\top_inst.deskew_buff_inst.col_input[40] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\top_inst.axis_out_inst.out_buff_data[103] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\top_inst.axis_out_inst.out_buff_data[53] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][5] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][11] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][17] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][0] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\top_inst.deskew_buff_inst.col_input[83] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][25] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][7] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\top_inst.skew_buff_inst.row[1].has_delay.shift_reg[0][5] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(_00963_),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\top_inst.deskew_buff_inst.col_input[41] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\top_inst.deskew_buff_inst.col_input[118] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][17] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\top_inst.deskew_buff_inst.col_input[84] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(_00059_),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][2] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][24] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][16] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\top_inst.deskew_buff_inst.col_input[81] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][5] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\top_inst.deskew_buff_inst.col_input[106] ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\top_inst.deskew_buff_inst.col_input[37] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][27] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][6] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\top_inst.deskew_buff_inst.col_input[74] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][4] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(_00906_),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][24] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][7] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\top_inst.axis_in_inst.inbuf_bus[11] ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\top_inst.axis_in_inst.inbuf_bus[0] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(_00974_),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][8] ),
    .X(net905));
 sky130_fd_sc_hd__buf_1 hold724 (.A(\top_inst.deskew_buff_inst.col_input[26] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\top_inst.deskew_buff_inst.col_input[19] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][21] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][8] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][26] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\top_inst.deskew_buff_inst.col_input[6] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[1][4] ),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][14] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][20] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(_00091_),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][9] ),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\top_inst.deskew_buff_inst.col_input[0] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\top_inst.axis_in_inst.inbuf_bus[19] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\top_inst.deskew_buff_inst.col_input[57] ),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\top_inst.axis_out_inst.out_buff_data[59] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\top_inst.deskew_buff_inst.col_input[69] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[17] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\top_inst.deskew_buff_inst.col_input[113] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\top_inst.deskew_buff_inst.col_input[73] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\top_inst.deskew_buff_inst.col_input[20] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][14] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\top_inst.axis_out_inst.out_buff_data[80] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[19] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][31] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[2][0] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(_00167_),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\top_inst.deskew_buff_inst.col_input[1] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][20] ),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\top_inst.deskew_buff_inst.col_input[23] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[1] ),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\top_inst.skew_buff_inst.row[3].has_delay.shift_reg[2][0] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(_00902_),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\top_inst.deskew_buff_inst.col_input[71] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[19] ),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(\top_inst.axis_out_inst.out_buff_data[68] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][12] ),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(\top_inst.axis_in_inst.inbuf_bus[25] ),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\top_inst.deskew_buff_inst.row[0].delayed_pass.shift_reg[0][15] ),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(\top_inst.deskew_buff_inst.row[2].delayed_pass.shift_reg[0][28] ),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\top_inst.axis_out_inst.out_buff_data[55] ),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[17] ),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[20] ),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[18] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[24] ),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[0] ),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\top_inst.axis_in_inst.inbuf_bus[2] ),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(_00976_),
    .X(net952));
 sky130_fd_sc_hd__buf_1 hold771 (.A(\top_inst.deskew_buff_inst.col_input[89] ),
    .X(net953));
 sky130_fd_sc_hd__buf_1 hold772 (.A(\top_inst.deskew_buff_inst.col_input[95] ),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\top_inst.axis_out_inst.out_buff_data[15] ),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[18] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[18] ),
    .X(net957));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold776 (.A(\top_inst.deskew_buff_inst.col_input[21] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[19] ),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[20] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[21] ),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[23] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[17] ),
    .X(net963));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold782 (.A(\top_inst.deskew_buff_inst.col_input[105] ),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\top_inst.axis_in_inst.inbuf_bus[12] ),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(\top_inst.deskew_buff_inst.col_input[51] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][16] ),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(\top_inst.deskew_buff_inst.col_input[17] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\top_inst.axis_in_inst.inbuf_bus[10] ),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][6] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\top_inst.axis_in_inst.inbuf_bus[15] ),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\top_inst.axis_out_inst.out_buff_data[31] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][26] ),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[13] ),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[23] ),
    .X(net975));
 sky130_fd_sc_hd__buf_1 hold794 (.A(\top_inst.deskew_buff_inst.col_input[25] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[1] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(\top_inst.axis_out_inst.out_buff_data[52] ),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\top_inst.axis_in_inst.inbuf_bus[3] ),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(_00977_),
    .X(net980));
 sky130_fd_sc_hd__buf_1 hold799 (.A(\top_inst.deskew_buff_inst.col_input[27] ),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[6] ),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\top_inst.axis_in_inst.inbuf_bus[1] ),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(_00975_),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[24] ),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(\top_inst.axis_in_inst.inbuf_bus[29] ),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\top_inst.axis_in_inst.inbuf_bus[24] ),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(\top_inst.axis_out_inst.out_buff_data[0] ),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[31] ),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[0] ),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\top_inst.axis_in_inst.inbuf_bus[17] ),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(\top_inst.axis_in_inst.inbuf_bus[9] ),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\top_inst.axis_out_inst.out_buff_data[99] ),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(\top_inst.axis_in_inst.inbuf_bus[18] ),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\top_inst.axis_in_inst.inbuf_bus[13] ),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[0] ),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\top_inst.deskew_buff_inst.col_input[59] ),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[14] ),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][10] ),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[1] ),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][1] ),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[20] ),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\top_inst.axis_in_inst.inbuf_bus[30] ),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[1] ),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[2] ),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(\top_inst.axis_in_inst.inbuf_bus[31] ),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\top_inst.axis_in_inst.inbuf_bus[21] ),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[13] ),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[23] ),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[10] ),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[13] ),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][11] ),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[8] ),
    .X(net1013));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold832 (.A(\top_inst.deskew_buff_inst.col_input[96] ),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\top_inst.axis_in_inst.inbuf_bus[23] ),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[9] ),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[0] ),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[21] ),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\top_inst.axis_in_inst.inbuf_bus[4] ),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(_00978_),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][12] ),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[17] ),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\top_inst.axis_out_inst.out_buff_data[63] ),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[9] ),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\top_inst.axis_out_inst.out_buff_data[58] ),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[1] ),
    .X(net1026));
 sky130_fd_sc_hd__buf_1 hold845 (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[1] ),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[27] ),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\top_inst.axis_in_inst.inbuf_bus[16] ),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[28] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[3] ),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[27] ),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[11] ),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(\top_inst.axis_in_inst.inbuf_bus[27] ),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[15] ),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[2] ),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\top_inst.axis_in_inst.inbuf_bus[22] ),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[11] ),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\top_inst.axis_in_inst.inbuf_bus[26] ),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[11] ),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[0] ),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[15] ),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\top_inst.axis_in_inst.inbuf_bus[28] ),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[0] ),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[1] ),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[21] ),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[23] ),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[3] ),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[13] ),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[21] ),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[25] ),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[11] ),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[4] ),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[13] ),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[15] ),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[2] ),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\top_inst.grid_inst.rows[2].cols[3].pe_inst.sum_output[25] ),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.weight_reg[7] ),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\top_inst.axis_out_inst.out_buff_data[61] ),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[1] ),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[9] ),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[14] ),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\top_inst.skew_buff_inst.row[0].output_reg[6] ),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[1] ),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[12] ),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[13] ),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[15] ),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(\top_inst.grid_inst.rows[1].cols[3].pe_inst.sum_output[0] ),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(_00532_),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[4] ),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\top_inst.grid_inst.rows[1].cols[1].pe_inst.sum_output[4] ),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[3] ),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[3] ),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(\top_inst.grid_inst.rows[0].cols[2].pe_inst.sum_output[15] ),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[0] ),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[25] ),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[0] ),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[0] ),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[2] ),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[16] ),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[4] ),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[17] ),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[10] ),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(\top_inst.grid_inst.rows[0].cols[0].pe_inst.sum_output[9] ),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\top_inst.grid_inst.rows[2].cols[2].pe_inst.sum_output[13] ),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(\top_inst.grid_inst.rows[1].cols[2].pe_inst.sum_output[9] ),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\top_inst.grid_inst.rows[0].cols[1].pe_inst.sum_output[2] ),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(\top_inst.grid_inst.rows[1].cols[0].pe_inst.sum_output[15] ),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\top_inst.grid_inst.rows[2].cols[1].pe_inst.sum_output[12] ),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(\top_inst.grid_inst.rows[0].cols[3].pe_inst.sum_output[12] ),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\top_inst.grid_inst.rows[2].cols[0].pe_inst.sum_output[12] ),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(\top_inst.deskew_buff_inst.col_input[11] ),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\top_inst.deskew_buff_inst.col_input[15] ),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(\top_inst.deskew_buff_inst.col_input[23] ),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\top_inst.deskew_buff_inst.col_input[21] ),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(\top_inst.deskew_buff_inst.col_input[17] ),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\top_inst.deskew_buff_inst.col_input[62] ),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(\top_inst.deskew_buff_inst.col_input[27] ),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\top_inst.deskew_buff_inst.col_input[25] ),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][10] ),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\top_inst.axis_out_inst.out_buff_data[58] ),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(\top_inst.deskew_buff_inst.col_input[63] ),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\top_inst.deskew_buff_inst.col_input[98] ),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][11] ),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[0][19] ),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(\top_inst.deskew_buff_inst.row[1].delayed_pass.shift_reg[1][12] ),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\top_inst.axis_out_inst.out_buff_data[99] ),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(\top_inst.axis_out_inst.out_buff_data[63] ),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\top_inst.axis_in_inst.inbuf_bus[21] ),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(\top_inst.axis_in_inst.inbuf_bus[23] ),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\top_inst.axis_in_inst.inbuf_bus[19] ),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(\top_inst.axis_in_inst.inbuf_bus[7] ),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\top_inst.axis_in_inst.inbuf_bus[31] ),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(\top_inst.axis_in_inst.inbuf_bus[27] ),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\top_inst.axis_in_inst.inbuf_bus[30] ),
    .X(net1115));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer6 (.A(_09892_),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(net1116),
    .X(net253));
 sky130_fd_sc_hd__buf_2 rebuffer47 (.A(_01464_),
    .X(net1116));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer70 (.A(_09560_),
    .X(net1117));
 sky130_fd_sc_hd__buf_2 rebuffer71 (.A(_09529_),
    .X(net1118));
 sky130_fd_sc_hd__buf_1 rebuffer72 (.A(_09191_),
    .X(net1119));
 sky130_fd_sc_hd__buf_2 rebuffer73 (.A(net1119),
    .X(net1120));
 sky130_fd_sc_hd__clkbuf_1 rebuffer74 (.A(_09559_),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer75 (.A(_07081_),
    .X(net1122));
 sky130_fd_sc_hd__clkbuf_1 rebuffer76 (.A(net1122),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer77 (.A(_07437_),
    .X(net1124));
 sky130_fd_sc_hd__clkbuf_2 rebuffer78 (.A(_07151_),
    .X(net1125));
 sky130_fd_sc_hd__clkbuf_1 rebuffer79 (.A(_01416_),
    .X(net1126));
endmodule
