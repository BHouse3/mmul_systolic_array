VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_hardened
  CLASS BLOCK ;
  FOREIGN top_hardened ;
  ORIGIN 0.000 0.000 ;
  SIZE 678.570 BY 689.290 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 677.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 677.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 677.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 677.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 677.520 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 673.220 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 673.220 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 673.220 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 489.570 673.220 491.170 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 642.750 673.220 644.350 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 677.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 677.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 677.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 677.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 677.520 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 673.220 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 673.220 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 673.220 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 673.220 487.870 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 639.450 673.220 641.050 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END clk
  PIN input_tdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 674.570 173.440 678.570 174.040 ;
    END
  END input_tdata[0]
  PIN input_tdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 105.440 678.570 106.040 ;
    END
  END input_tdata[10]
  PIN input_tdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END input_tdata[11]
  PIN input_tdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END input_tdata[12]
  PIN input_tdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 674.570 629.040 678.570 629.640 ;
    END
  END input_tdata[13]
  PIN input_tdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 674.570 544.040 678.570 544.640 ;
    END
  END input_tdata[14]
  PIN input_tdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END input_tdata[15]
  PIN input_tdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 524.950 685.290 525.230 689.290 ;
    END
  END input_tdata[16]
  PIN input_tdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 383.270 685.290 383.550 689.290 ;
    END
  END input_tdata[17]
  PIN input_tdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END input_tdata[18]
  PIN input_tdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 74.840 678.570 75.440 ;
    END
  END input_tdata[19]
  PIN input_tdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 589.350 685.290 589.630 689.290 ;
    END
  END input_tdata[1]
  PIN input_tdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END input_tdata[20]
  PIN input_tdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 674.570 561.040 678.570 561.640 ;
    END
  END input_tdata[21]
  PIN input_tdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END input_tdata[22]
  PIN input_tdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END input_tdata[23]
  PIN input_tdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 96.690 685.290 96.970 689.290 ;
    END
  END input_tdata[24]
  PIN input_tdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END input_tdata[25]
  PIN input_tdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END input_tdata[26]
  PIN input_tdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 351.070 685.290 351.350 689.290 ;
    END
  END input_tdata[27]
  PIN input_tdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 190.070 685.290 190.350 689.290 ;
    END
  END input_tdata[28]
  PIN input_tdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END input_tdata[29]
  PIN input_tdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END input_tdata[2]
  PIN input_tdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 674.570 40.840 678.570 41.440 ;
    END
  END input_tdata[30]
  PIN input_tdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END input_tdata[31]
  PIN input_tdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 447.670 685.290 447.950 689.290 ;
    END
  END input_tdata[3]
  PIN input_tdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END input_tdata[4]
  PIN input_tdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 674.570 343.440 678.570 344.040 ;
    END
  END input_tdata[5]
  PIN input_tdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END input_tdata[6]
  PIN input_tdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 674.570 394.440 678.570 395.040 ;
    END
  END input_tdata[7]
  PIN input_tdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 286.670 685.290 286.950 689.290 ;
    END
  END input_tdata[8]
  PIN input_tdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END input_tdata[9]
  PIN input_tready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END input_tready
  PIN input_tvalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 621.550 685.290 621.830 689.290 ;
    END
  END input_tvalid
  PIN load_weight
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 302.770 685.290 303.050 689.290 ;
    END
  END load_weight
  PIN output_tdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END output_tdata[0]
  PIN output_tdata[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 206.170 685.290 206.450 689.290 ;
    END
  END output_tdata[100]
  PIN output_tdata[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END output_tdata[101]
  PIN output_tdata[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END output_tdata[102]
  PIN output_tdata[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 173.970 685.290 174.250 689.290 ;
    END
  END output_tdata[103]
  PIN output_tdata[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 674.570 309.440 678.570 310.040 ;
    END
  END output_tdata[104]
  PIN output_tdata[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 222.270 685.290 222.550 689.290 ;
    END
  END output_tdata[105]
  PIN output_tdata[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 527.040 678.570 527.640 ;
    END
  END output_tdata[106]
  PIN output_tdata[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 428.440 678.570 429.040 ;
    END
  END output_tdata[107]
  PIN output_tdata[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END output_tdata[108]
  PIN output_tdata[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END output_tdata[109]
  PIN output_tdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END output_tdata[10]
  PIN output_tdata[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END output_tdata[110]
  PIN output_tdata[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 674.570 88.440 678.570 89.040 ;
    END
  END output_tdata[111]
  PIN output_tdata[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END output_tdata[112]
  PIN output_tdata[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END output_tdata[113]
  PIN output_tdata[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 637.650 685.290 637.930 689.290 ;
    END
  END output_tdata[114]
  PIN output_tdata[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END output_tdata[115]
  PIN output_tdata[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END output_tdata[116]
  PIN output_tdata[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END output_tdata[117]
  PIN output_tdata[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 653.750 685.290 654.030 689.290 ;
    END
  END output_tdata[118]
  PIN output_tdata[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 669.850 685.290 670.130 689.290 ;
    END
  END output_tdata[119]
  PIN output_tdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 64.490 685.290 64.770 689.290 ;
    END
  END output_tdata[11]
  PIN output_tdata[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 318.870 685.290 319.150 689.290 ;
    END
  END output_tdata[120]
  PIN output_tdata[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 80.590 685.290 80.870 689.290 ;
    END
  END output_tdata[121]
  PIN output_tdata[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END output_tdata[122]
  PIN output_tdata[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 674.570 275.440 678.570 276.040 ;
    END
  END output_tdata[123]
  PIN output_tdata[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 431.570 685.290 431.850 689.290 ;
    END
  END output_tdata[124]
  PIN output_tdata[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 16.190 685.290 16.470 689.290 ;
    END
  END output_tdata[125]
  PIN output_tdata[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 463.770 685.290 464.050 689.290 ;
    END
  END output_tdata[126]
  PIN output_tdata[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 360.440 678.570 361.040 ;
    END
  END output_tdata[127]
  PIN output_tdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 663.040 678.570 663.640 ;
    END
  END output_tdata[12]
  PIN output_tdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END output_tdata[13]
  PIN output_tdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 605.450 685.290 605.730 689.290 ;
    END
  END output_tdata[14]
  PIN output_tdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END output_tdata[15]
  PIN output_tdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END output_tdata[16]
  PIN output_tdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END output_tdata[17]
  PIN output_tdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 612.040 678.570 612.640 ;
    END
  END output_tdata[18]
  PIN output_tdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END output_tdata[19]
  PIN output_tdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 241.440 678.570 242.040 ;
    END
  END output_tdata[1]
  PIN output_tdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 270.570 685.290 270.850 689.290 ;
    END
  END output_tdata[20]
  PIN output_tdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END output_tdata[21]
  PIN output_tdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END output_tdata[22]
  PIN output_tdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END output_tdata[23]
  PIN output_tdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 674.570 510.040 678.570 510.640 ;
    END
  END output_tdata[24]
  PIN output_tdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END output_tdata[25]
  PIN output_tdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END output_tdata[26]
  PIN output_tdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END output_tdata[27]
  PIN output_tdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END output_tdata[28]
  PIN output_tdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 674.570 156.440 678.570 157.040 ;
    END
  END output_tdata[29]
  PIN output_tdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 141.770 685.290 142.050 689.290 ;
    END
  END output_tdata[2]
  PIN output_tdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 292.440 678.570 293.040 ;
    END
  END output_tdata[30]
  PIN output_tdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END output_tdata[31]
  PIN output_tdata[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 157.870 685.290 158.150 689.290 ;
    END
  END output_tdata[32]
  PIN output_tdata[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END output_tdata[33]
  PIN output_tdata[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END output_tdata[34]
  PIN output_tdata[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END output_tdata[35]
  PIN output_tdata[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 399.370 685.290 399.650 689.290 ;
    END
  END output_tdata[36]
  PIN output_tdata[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END output_tdata[37]
  PIN output_tdata[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END output_tdata[38]
  PIN output_tdata[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 595.040 678.570 595.640 ;
    END
  END output_tdata[39]
  PIN output_tdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 207.440 678.570 208.040 ;
    END
  END output_tdata[3]
  PIN output_tdata[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 415.470 685.290 415.750 689.290 ;
    END
  END output_tdata[40]
  PIN output_tdata[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 508.850 685.290 509.130 689.290 ;
    END
  END output_tdata[41]
  PIN output_tdata[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END output_tdata[42]
  PIN output_tdata[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END output_tdata[43]
  PIN output_tdata[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END output_tdata[44]
  PIN output_tdata[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 57.840 678.570 58.440 ;
    END
  END output_tdata[45]
  PIN output_tdata[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 32.290 685.290 32.570 689.290 ;
    END
  END output_tdata[46]
  PIN output_tdata[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 493.040 678.570 493.640 ;
    END
  END output_tdata[47]
  PIN output_tdata[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 238.370 685.290 238.650 689.290 ;
    END
  END output_tdata[48]
  PIN output_tdata[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 541.050 685.290 541.330 689.290 ;
    END
  END output_tdata[49]
  PIN output_tdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 48.390 685.290 48.670 689.290 ;
    END
  END output_tdata[4]
  PIN output_tdata[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 139.440 678.570 140.040 ;
    END
  END output_tdata[50]
  PIN output_tdata[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 674.570 377.440 678.570 378.040 ;
    END
  END output_tdata[51]
  PIN output_tdata[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 254.470 685.290 254.750 689.290 ;
    END
  END output_tdata[52]
  PIN output_tdata[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 258.440 678.570 259.040 ;
    END
  END output_tdata[53]
  PIN output_tdata[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 674.570 6.840 678.570 7.440 ;
    END
  END output_tdata[54]
  PIN output_tdata[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END output_tdata[55]
  PIN output_tdata[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 479.440 678.570 480.040 ;
    END
  END output_tdata[56]
  PIN output_tdata[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 557.150 685.290 557.430 689.290 ;
    END
  END output_tdata[57]
  PIN output_tdata[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END output_tdata[58]
  PIN output_tdata[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 190.440 678.570 191.040 ;
    END
  END output_tdata[59]
  PIN output_tdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END output_tdata[5]
  PIN output_tdata[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 23.840 678.570 24.440 ;
    END
  END output_tdata[60]
  PIN output_tdata[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 125.670 685.290 125.950 689.290 ;
    END
  END output_tdata[61]
  PIN output_tdata[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END output_tdata[62]
  PIN output_tdata[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END output_tdata[63]
  PIN output_tdata[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END output_tdata[64]
  PIN output_tdata[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END output_tdata[65]
  PIN output_tdata[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 674.570 578.040 678.570 578.640 ;
    END
  END output_tdata[66]
  PIN output_tdata[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 411.440 678.570 412.040 ;
    END
  END output_tdata[67]
  PIN output_tdata[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END output_tdata[68]
  PIN output_tdata[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END output_tdata[69]
  PIN output_tdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 224.440 678.570 225.040 ;
    END
  END output_tdata[6]
  PIN output_tdata[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END output_tdata[70]
  PIN output_tdata[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 445.440 678.570 446.040 ;
    END
  END output_tdata[71]
  PIN output_tdata[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 646.040 678.570 646.640 ;
    END
  END output_tdata[72]
  PIN output_tdata[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END output_tdata[73]
  PIN output_tdata[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 674.570 680.040 678.570 680.640 ;
    END
  END output_tdata[74]
  PIN output_tdata[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END output_tdata[75]
  PIN output_tdata[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END output_tdata[76]
  PIN output_tdata[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END output_tdata[77]
  PIN output_tdata[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END output_tdata[78]
  PIN output_tdata[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END output_tdata[79]
  PIN output_tdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END output_tdata[7]
  PIN output_tdata[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END output_tdata[80]
  PIN output_tdata[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 367.170 685.290 367.450 689.290 ;
    END
  END output_tdata[81]
  PIN output_tdata[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END output_tdata[82]
  PIN output_tdata[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END output_tdata[83]
  PIN output_tdata[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END output_tdata[84]
  PIN output_tdata[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END output_tdata[85]
  PIN output_tdata[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 334.970 685.290 335.250 689.290 ;
    END
  END output_tdata[86]
  PIN output_tdata[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END output_tdata[87]
  PIN output_tdata[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 573.250 685.290 573.530 689.290 ;
    END
  END output_tdata[88]
  PIN output_tdata[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 122.440 678.570 123.040 ;
    END
  END output_tdata[89]
  PIN output_tdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END output_tdata[8]
  PIN output_tdata[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END output_tdata[90]
  PIN output_tdata[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END output_tdata[91]
  PIN output_tdata[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END output_tdata[92]
  PIN output_tdata[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END output_tdata[93]
  PIN output_tdata[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 674.570 462.440 678.570 463.040 ;
    END
  END output_tdata[94]
  PIN output_tdata[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END output_tdata[95]
  PIN output_tdata[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 492.750 685.290 493.030 689.290 ;
    END
  END output_tdata[96]
  PIN output_tdata[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 479.870 685.290 480.150 689.290 ;
    END
  END output_tdata[97]
  PIN output_tdata[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 685.290 0.370 689.290 ;
    END
  END output_tdata[98]
  PIN output_tdata[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 109.570 685.290 109.850 689.290 ;
    END
  END output_tdata[99]
  PIN output_tdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END output_tdata[9]
  PIN output_tready
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END output_tready
  PIN output_tvalid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END output_tvalid
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 674.570 326.440 678.570 327.040 ;
    END
  END reset
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 672.980 677.365 ;
      LAYER met1 ;
        RECT 0.070 9.560 673.830 677.520 ;
      LAYER met2 ;
        RECT 0.650 685.010 15.910 685.850 ;
        RECT 16.750 685.010 32.010 685.850 ;
        RECT 32.850 685.010 48.110 685.850 ;
        RECT 48.950 685.010 64.210 685.850 ;
        RECT 65.050 685.010 80.310 685.850 ;
        RECT 81.150 685.010 96.410 685.850 ;
        RECT 97.250 685.010 109.290 685.850 ;
        RECT 110.130 685.010 125.390 685.850 ;
        RECT 126.230 685.010 141.490 685.850 ;
        RECT 142.330 685.010 157.590 685.850 ;
        RECT 158.430 685.010 173.690 685.850 ;
        RECT 174.530 685.010 189.790 685.850 ;
        RECT 190.630 685.010 205.890 685.850 ;
        RECT 206.730 685.010 221.990 685.850 ;
        RECT 222.830 685.010 238.090 685.850 ;
        RECT 238.930 685.010 254.190 685.850 ;
        RECT 255.030 685.010 270.290 685.850 ;
        RECT 271.130 685.010 286.390 685.850 ;
        RECT 287.230 685.010 302.490 685.850 ;
        RECT 303.330 685.010 318.590 685.850 ;
        RECT 319.430 685.010 334.690 685.850 ;
        RECT 335.530 685.010 350.790 685.850 ;
        RECT 351.630 685.010 366.890 685.850 ;
        RECT 367.730 685.010 382.990 685.850 ;
        RECT 383.830 685.010 399.090 685.850 ;
        RECT 399.930 685.010 415.190 685.850 ;
        RECT 416.030 685.010 431.290 685.850 ;
        RECT 432.130 685.010 447.390 685.850 ;
        RECT 448.230 685.010 463.490 685.850 ;
        RECT 464.330 685.010 479.590 685.850 ;
        RECT 480.430 685.010 492.470 685.850 ;
        RECT 493.310 685.010 508.570 685.850 ;
        RECT 509.410 685.010 524.670 685.850 ;
        RECT 525.510 685.010 540.770 685.850 ;
        RECT 541.610 685.010 556.870 685.850 ;
        RECT 557.710 685.010 572.970 685.850 ;
        RECT 573.810 685.010 589.070 685.850 ;
        RECT 589.910 685.010 605.170 685.850 ;
        RECT 606.010 685.010 621.270 685.850 ;
        RECT 622.110 685.010 637.370 685.850 ;
        RECT 638.210 685.010 653.470 685.850 ;
        RECT 654.310 685.010 669.570 685.850 ;
        RECT 670.410 685.010 673.810 685.850 ;
        RECT 0.100 4.280 673.810 685.010 ;
        RECT 0.650 3.670 12.690 4.280 ;
        RECT 13.530 3.670 28.790 4.280 ;
        RECT 29.630 3.670 44.890 4.280 ;
        RECT 45.730 3.670 60.990 4.280 ;
        RECT 61.830 3.670 77.090 4.280 ;
        RECT 77.930 3.670 93.190 4.280 ;
        RECT 94.030 3.670 109.290 4.280 ;
        RECT 110.130 3.670 125.390 4.280 ;
        RECT 126.230 3.670 141.490 4.280 ;
        RECT 142.330 3.670 157.590 4.280 ;
        RECT 158.430 3.670 173.690 4.280 ;
        RECT 174.530 3.670 189.790 4.280 ;
        RECT 190.630 3.670 205.890 4.280 ;
        RECT 206.730 3.670 221.990 4.280 ;
        RECT 222.830 3.670 238.090 4.280 ;
        RECT 238.930 3.670 254.190 4.280 ;
        RECT 255.030 3.670 270.290 4.280 ;
        RECT 271.130 3.670 286.390 4.280 ;
        RECT 287.230 3.670 302.490 4.280 ;
        RECT 303.330 3.670 318.590 4.280 ;
        RECT 319.430 3.670 334.690 4.280 ;
        RECT 335.530 3.670 350.790 4.280 ;
        RECT 351.630 3.670 366.890 4.280 ;
        RECT 367.730 3.670 379.770 4.280 ;
        RECT 380.610 3.670 395.870 4.280 ;
        RECT 396.710 3.670 411.970 4.280 ;
        RECT 412.810 3.670 428.070 4.280 ;
        RECT 428.910 3.670 444.170 4.280 ;
        RECT 445.010 3.670 460.270 4.280 ;
        RECT 461.110 3.670 476.370 4.280 ;
        RECT 477.210 3.670 492.470 4.280 ;
        RECT 493.310 3.670 508.570 4.280 ;
        RECT 509.410 3.670 524.670 4.280 ;
        RECT 525.510 3.670 540.770 4.280 ;
        RECT 541.610 3.670 556.870 4.280 ;
        RECT 557.710 3.670 572.970 4.280 ;
        RECT 573.810 3.670 589.070 4.280 ;
        RECT 589.910 3.670 605.170 4.280 ;
        RECT 606.010 3.670 621.270 4.280 ;
        RECT 622.110 3.670 637.370 4.280 ;
        RECT 638.210 3.670 653.470 4.280 ;
        RECT 654.310 3.670 669.570 4.280 ;
        RECT 670.410 3.670 673.810 4.280 ;
      LAYER met3 ;
        RECT 3.990 679.640 674.170 680.505 ;
        RECT 3.990 674.240 674.570 679.640 ;
        RECT 4.400 672.840 674.570 674.240 ;
        RECT 3.990 664.040 674.570 672.840 ;
        RECT 3.990 662.640 674.170 664.040 ;
        RECT 3.990 657.240 674.570 662.640 ;
        RECT 4.400 655.840 674.570 657.240 ;
        RECT 3.990 647.040 674.570 655.840 ;
        RECT 3.990 645.640 674.170 647.040 ;
        RECT 3.990 640.240 674.570 645.640 ;
        RECT 4.400 638.840 674.570 640.240 ;
        RECT 3.990 630.040 674.570 638.840 ;
        RECT 3.990 628.640 674.170 630.040 ;
        RECT 3.990 623.240 674.570 628.640 ;
        RECT 4.400 621.840 674.570 623.240 ;
        RECT 3.990 613.040 674.570 621.840 ;
        RECT 3.990 611.640 674.170 613.040 ;
        RECT 3.990 606.240 674.570 611.640 ;
        RECT 4.400 604.840 674.570 606.240 ;
        RECT 3.990 596.040 674.570 604.840 ;
        RECT 3.990 594.640 674.170 596.040 ;
        RECT 3.990 589.240 674.570 594.640 ;
        RECT 4.400 587.840 674.570 589.240 ;
        RECT 3.990 579.040 674.570 587.840 ;
        RECT 3.990 577.640 674.170 579.040 ;
        RECT 3.990 572.240 674.570 577.640 ;
        RECT 4.400 570.840 674.570 572.240 ;
        RECT 3.990 562.040 674.570 570.840 ;
        RECT 3.990 560.640 674.170 562.040 ;
        RECT 3.990 555.240 674.570 560.640 ;
        RECT 4.400 553.840 674.570 555.240 ;
        RECT 3.990 545.040 674.570 553.840 ;
        RECT 3.990 543.640 674.170 545.040 ;
        RECT 3.990 538.240 674.570 543.640 ;
        RECT 4.400 536.840 674.570 538.240 ;
        RECT 3.990 528.040 674.570 536.840 ;
        RECT 3.990 526.640 674.170 528.040 ;
        RECT 3.990 521.240 674.570 526.640 ;
        RECT 4.400 519.840 674.570 521.240 ;
        RECT 3.990 511.040 674.570 519.840 ;
        RECT 3.990 509.640 674.170 511.040 ;
        RECT 3.990 504.240 674.570 509.640 ;
        RECT 4.400 502.840 674.570 504.240 ;
        RECT 3.990 494.040 674.570 502.840 ;
        RECT 3.990 492.640 674.170 494.040 ;
        RECT 3.990 487.240 674.570 492.640 ;
        RECT 4.400 485.840 674.570 487.240 ;
        RECT 3.990 480.440 674.570 485.840 ;
        RECT 3.990 479.040 674.170 480.440 ;
        RECT 3.990 470.240 674.570 479.040 ;
        RECT 4.400 468.840 674.570 470.240 ;
        RECT 3.990 463.440 674.570 468.840 ;
        RECT 3.990 462.040 674.170 463.440 ;
        RECT 3.990 453.240 674.570 462.040 ;
        RECT 4.400 451.840 674.570 453.240 ;
        RECT 3.990 446.440 674.570 451.840 ;
        RECT 3.990 445.040 674.170 446.440 ;
        RECT 3.990 436.240 674.570 445.040 ;
        RECT 4.400 434.840 674.570 436.240 ;
        RECT 3.990 429.440 674.570 434.840 ;
        RECT 3.990 428.040 674.170 429.440 ;
        RECT 3.990 419.240 674.570 428.040 ;
        RECT 4.400 417.840 674.570 419.240 ;
        RECT 3.990 412.440 674.570 417.840 ;
        RECT 3.990 411.040 674.170 412.440 ;
        RECT 3.990 402.240 674.570 411.040 ;
        RECT 4.400 400.840 674.570 402.240 ;
        RECT 3.990 395.440 674.570 400.840 ;
        RECT 3.990 394.040 674.170 395.440 ;
        RECT 3.990 388.640 674.570 394.040 ;
        RECT 4.400 387.240 674.570 388.640 ;
        RECT 3.990 378.440 674.570 387.240 ;
        RECT 3.990 377.040 674.170 378.440 ;
        RECT 3.990 371.640 674.570 377.040 ;
        RECT 4.400 370.240 674.570 371.640 ;
        RECT 3.990 361.440 674.570 370.240 ;
        RECT 3.990 360.040 674.170 361.440 ;
        RECT 3.990 354.640 674.570 360.040 ;
        RECT 4.400 353.240 674.570 354.640 ;
        RECT 3.990 344.440 674.570 353.240 ;
        RECT 3.990 343.040 674.170 344.440 ;
        RECT 3.990 337.640 674.570 343.040 ;
        RECT 4.400 336.240 674.570 337.640 ;
        RECT 3.990 327.440 674.570 336.240 ;
        RECT 3.990 326.040 674.170 327.440 ;
        RECT 3.990 320.640 674.570 326.040 ;
        RECT 4.400 319.240 674.570 320.640 ;
        RECT 3.990 310.440 674.570 319.240 ;
        RECT 3.990 309.040 674.170 310.440 ;
        RECT 3.990 303.640 674.570 309.040 ;
        RECT 4.400 302.240 674.570 303.640 ;
        RECT 3.990 293.440 674.570 302.240 ;
        RECT 3.990 292.040 674.170 293.440 ;
        RECT 3.990 286.640 674.570 292.040 ;
        RECT 4.400 285.240 674.570 286.640 ;
        RECT 3.990 276.440 674.570 285.240 ;
        RECT 3.990 275.040 674.170 276.440 ;
        RECT 3.990 269.640 674.570 275.040 ;
        RECT 4.400 268.240 674.570 269.640 ;
        RECT 3.990 259.440 674.570 268.240 ;
        RECT 3.990 258.040 674.170 259.440 ;
        RECT 3.990 252.640 674.570 258.040 ;
        RECT 4.400 251.240 674.570 252.640 ;
        RECT 3.990 242.440 674.570 251.240 ;
        RECT 3.990 241.040 674.170 242.440 ;
        RECT 3.990 235.640 674.570 241.040 ;
        RECT 4.400 234.240 674.570 235.640 ;
        RECT 3.990 225.440 674.570 234.240 ;
        RECT 3.990 224.040 674.170 225.440 ;
        RECT 3.990 218.640 674.570 224.040 ;
        RECT 4.400 217.240 674.570 218.640 ;
        RECT 3.990 208.440 674.570 217.240 ;
        RECT 3.990 207.040 674.170 208.440 ;
        RECT 3.990 201.640 674.570 207.040 ;
        RECT 4.400 200.240 674.570 201.640 ;
        RECT 3.990 191.440 674.570 200.240 ;
        RECT 3.990 190.040 674.170 191.440 ;
        RECT 3.990 184.640 674.570 190.040 ;
        RECT 4.400 183.240 674.570 184.640 ;
        RECT 3.990 174.440 674.570 183.240 ;
        RECT 3.990 173.040 674.170 174.440 ;
        RECT 3.990 167.640 674.570 173.040 ;
        RECT 4.400 166.240 674.570 167.640 ;
        RECT 3.990 157.440 674.570 166.240 ;
        RECT 3.990 156.040 674.170 157.440 ;
        RECT 3.990 150.640 674.570 156.040 ;
        RECT 4.400 149.240 674.570 150.640 ;
        RECT 3.990 140.440 674.570 149.240 ;
        RECT 3.990 139.040 674.170 140.440 ;
        RECT 3.990 133.640 674.570 139.040 ;
        RECT 4.400 132.240 674.570 133.640 ;
        RECT 3.990 123.440 674.570 132.240 ;
        RECT 3.990 122.040 674.170 123.440 ;
        RECT 3.990 116.640 674.570 122.040 ;
        RECT 4.400 115.240 674.570 116.640 ;
        RECT 3.990 106.440 674.570 115.240 ;
        RECT 3.990 105.040 674.170 106.440 ;
        RECT 3.990 99.640 674.570 105.040 ;
        RECT 4.400 98.240 674.570 99.640 ;
        RECT 3.990 89.440 674.570 98.240 ;
        RECT 3.990 88.040 674.170 89.440 ;
        RECT 3.990 82.640 674.570 88.040 ;
        RECT 4.400 81.240 674.570 82.640 ;
        RECT 3.990 75.840 674.570 81.240 ;
        RECT 3.990 74.440 674.170 75.840 ;
        RECT 3.990 65.640 674.570 74.440 ;
        RECT 4.400 64.240 674.570 65.640 ;
        RECT 3.990 58.840 674.570 64.240 ;
        RECT 3.990 57.440 674.170 58.840 ;
        RECT 3.990 48.640 674.570 57.440 ;
        RECT 4.400 47.240 674.570 48.640 ;
        RECT 3.990 41.840 674.570 47.240 ;
        RECT 3.990 40.440 674.170 41.840 ;
        RECT 3.990 31.640 674.570 40.440 ;
        RECT 4.400 30.240 674.570 31.640 ;
        RECT 3.990 24.840 674.570 30.240 ;
        RECT 3.990 23.440 674.170 24.840 ;
        RECT 3.990 14.640 674.570 23.440 ;
        RECT 4.400 13.240 674.570 14.640 ;
        RECT 3.990 7.840 674.570 13.240 ;
        RECT 3.990 6.975 674.170 7.840 ;
      LAYER met4 ;
        RECT 16.855 11.735 20.640 675.745 ;
        RECT 23.040 11.735 23.940 675.745 ;
        RECT 26.340 11.735 174.240 675.745 ;
        RECT 176.640 11.735 177.540 675.745 ;
        RECT 179.940 11.735 327.840 675.745 ;
        RECT 330.240 11.735 331.140 675.745 ;
        RECT 333.540 11.735 481.440 675.745 ;
        RECT 483.840 11.735 484.740 675.745 ;
        RECT 487.140 11.735 635.040 675.745 ;
        RECT 637.440 11.735 638.340 675.745 ;
        RECT 640.740 11.735 642.785 675.745 ;
  END
END top_hardened
END LIBRARY

